`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Yankai Wang
// 
// Create Date: 2025/05/10 20:02:30
// Design Name: polar_code
// Module Name: Sorter
// Project Name: polar_code
// Target Devices: zcu106
// Tool Versions: 2023.2
// Description: 
//   L为2的排序器
//   排序算法采用简化冒泡排序算法，利用PM特性：
//   PM_{2l} < PM_{2l+1}
//   PM_{2l} < PM_{2l+2}
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//   
//////////////////////////////////////////////////////////////////////////////////


module Sorter2(
    PM_in,
    PM_out
);

/*******************************************************************************/
/*                              Parameter                                      */
/*******************************************************************************/
parameter  PM_WIDTH    = 8;
parameter  INDEX_WIDTH = 2;
localparam L           = 2;
/*******************************************************************************/
/*                              IO Direction                                   */
/*******************************************************************************/
input  [PM_WIDTH*2*L-1:0]               PM_in;
output [(PM_WIDTH+INDEX_WIDTH)*L-1:0]   PM_out;
/*******************************************************************************/
/*                              Signal Declaration                             */
/*******************************************************************************/
// 第零阶段
wire [PM_WIDTH-1:0] m0_0;
wire [PM_WIDTH-1:0] m1_0;
wire [PM_WIDTH-1:0] m2_0;
wire [PM_WIDTH-1:0] m3_0;

// 第一阶段
wire [PM_WIDTH+INDEX_WIDTH-1:0] m0_1;
wire [PM_WIDTH+INDEX_WIDTH-1:0] m1_1;
wire [PM_WIDTH+INDEX_WIDTH-1:0] m2_1;
wire [PM_WIDTH+INDEX_WIDTH-1:0] m3_1;
/*******************************************************************************/
/*                              Instance                                       */
/*******************************************************************************/
/*******************************************************************************/
/*                              Logic                                          */
/*******************************************************************************/
assign {m0_0, m1_0, m2_0, m3_0} = PM_in;
assign PM_out = {m0_1, m1_1};

// 第一阶段
assign m0_1 = {2'd0, m0_0};
CAS #(.PM_WIDTH(PM_WIDTH), .INDEX_WIDTH(INDEX_WIDTH)) CAS_11 (.Din0({2'd1, m1_0}), .Din1({2'd2, m2_0}), .Dout0(m1_1), .Dout1(m2_1));
assign m3_1 = {2'd3, m3_0};
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/04/05 16:57:45
// Design Name: 
// Module Name: stage_1_xor_unit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`include "defines.v"

module stage_1_xor_unit(
    input [`STAGE1_INPUT_WIDTH-1 : 0] i_stage_1_comp_in,  //compute input
    output [`STAGE1_OUTPUT_WIDTH-1 : 0] o_stage_1_comp_out //compute output
    );

assign o_stage_1_comp_out[0]=i_stage_1_comp_in[0];
assign o_stage_1_comp_out[1]=i_stage_1_comp_in[0];
assign o_stage_1_comp_out[2]=i_stage_1_comp_in[0];
assign o_stage_1_comp_out[3]=i_stage_1_comp_in[0];
assign o_stage_1_comp_out[4]=i_stage_1_comp_in[1];
assign o_stage_1_comp_out[5]=i_stage_1_comp_in[1];
assign o_stage_1_comp_out[6]=i_stage_1_comp_in[1];
assign o_stage_1_comp_out[7]=i_stage_1_comp_in[1];
assign o_stage_1_comp_out[8]=i_stage_1_comp_in[2];
assign o_stage_1_comp_out[9]=i_stage_1_comp_in[2];
assign o_stage_1_comp_out[10]=i_stage_1_comp_in[2];
assign o_stage_1_comp_out[11]=i_stage_1_comp_in[2];
assign o_stage_1_comp_out[12]=i_stage_1_comp_in[3];
assign o_stage_1_comp_out[13]=i_stage_1_comp_in[3];
assign o_stage_1_comp_out[14]=i_stage_1_comp_in[3];
assign o_stage_1_comp_out[15]=i_stage_1_comp_in[3];
assign o_stage_1_comp_out[16]=i_stage_1_comp_in[4]^i_stage_1_comp_in[5]^i_stage_1_comp_in[6];
assign o_stage_1_comp_out[17]=i_stage_1_comp_in[4]^i_stage_1_comp_in[6];
assign o_stage_1_comp_out[18]=i_stage_1_comp_in[5]^i_stage_1_comp_in[6];
assign o_stage_1_comp_out[19]=i_stage_1_comp_in[6];
assign o_stage_1_comp_out[20]=i_stage_1_comp_in[7];
assign o_stage_1_comp_out[21]=i_stage_1_comp_in[7];
assign o_stage_1_comp_out[22]=i_stage_1_comp_in[7];
assign o_stage_1_comp_out[23]=i_stage_1_comp_in[7];
assign o_stage_1_comp_out[24]=i_stage_1_comp_in[8];
assign o_stage_1_comp_out[25]=i_stage_1_comp_in[8];
assign o_stage_1_comp_out[26]=i_stage_1_comp_in[8];
assign o_stage_1_comp_out[27]=i_stage_1_comp_in[8];
assign o_stage_1_comp_out[28]=i_stage_1_comp_in[9];
assign o_stage_1_comp_out[29]=i_stage_1_comp_in[9];
assign o_stage_1_comp_out[30]=i_stage_1_comp_in[9];
assign o_stage_1_comp_out[31]=i_stage_1_comp_in[9];
assign o_stage_1_comp_out[32]=i_stage_1_comp_in[10];
assign o_stage_1_comp_out[33]=i_stage_1_comp_in[10];
assign o_stage_1_comp_out[34]=i_stage_1_comp_in[10];
assign o_stage_1_comp_out[35]=i_stage_1_comp_in[10];
assign o_stage_1_comp_out[36]=i_stage_1_comp_in[11]^i_stage_1_comp_in[12]^i_stage_1_comp_in[13];
assign o_stage_1_comp_out[37]=i_stage_1_comp_in[11]^i_stage_1_comp_in[13];
assign o_stage_1_comp_out[38]=i_stage_1_comp_in[12]^i_stage_1_comp_in[13];
assign o_stage_1_comp_out[39]=i_stage_1_comp_in[13];
assign o_stage_1_comp_out[40]=i_stage_1_comp_in[14]^i_stage_1_comp_in[15]^i_stage_1_comp_in[16]^i_stage_1_comp_in[17];
assign o_stage_1_comp_out[41]=i_stage_1_comp_in[15]^i_stage_1_comp_in[17];
assign o_stage_1_comp_out[42]=i_stage_1_comp_in[16]^i_stage_1_comp_in[17];
assign o_stage_1_comp_out[43]=i_stage_1_comp_in[17];
assign o_stage_1_comp_out[44]=i_stage_1_comp_in[18]^i_stage_1_comp_in[19];
assign o_stage_1_comp_out[45]=i_stage_1_comp_in[19];
assign o_stage_1_comp_out[46]=i_stage_1_comp_in[18]^i_stage_1_comp_in[19];
assign o_stage_1_comp_out[47]=i_stage_1_comp_in[19];
assign o_stage_1_comp_out[48]=i_stage_1_comp_in[20]^i_stage_1_comp_in[21];
assign o_stage_1_comp_out[49]=i_stage_1_comp_in[21];
assign o_stage_1_comp_out[50]=i_stage_1_comp_in[20]^i_stage_1_comp_in[21];
assign o_stage_1_comp_out[51]=i_stage_1_comp_in[21];
assign o_stage_1_comp_out[52]=i_stage_1_comp_in[22];
assign o_stage_1_comp_out[53]=i_stage_1_comp_in[22];
assign o_stage_1_comp_out[54]=i_stage_1_comp_in[22];
assign o_stage_1_comp_out[55]=i_stage_1_comp_in[22];
assign o_stage_1_comp_out[56]=i_stage_1_comp_in[23]^i_stage_1_comp_in[24]^i_stage_1_comp_in[25];
assign o_stage_1_comp_out[57]=i_stage_1_comp_in[23]^i_stage_1_comp_in[25];
assign o_stage_1_comp_out[58]=i_stage_1_comp_in[24]^i_stage_1_comp_in[25];
assign o_stage_1_comp_out[59]=i_stage_1_comp_in[25];
assign o_stage_1_comp_out[60]=i_stage_1_comp_in[26]^i_stage_1_comp_in[27]^i_stage_1_comp_in[28];
assign o_stage_1_comp_out[61]=i_stage_1_comp_in[26]^i_stage_1_comp_in[28];
assign o_stage_1_comp_out[62]=i_stage_1_comp_in[27]^i_stage_1_comp_in[28];
assign o_stage_1_comp_out[63]=i_stage_1_comp_in[28];
assign o_stage_1_comp_out[64]=i_stage_1_comp_in[29]^i_stage_1_comp_in[30]^i_stage_1_comp_in[31]^i_stage_1_comp_in[32];
assign o_stage_1_comp_out[65]=i_stage_1_comp_in[30]^i_stage_1_comp_in[32];
assign o_stage_1_comp_out[66]=i_stage_1_comp_in[31]^i_stage_1_comp_in[32];
assign o_stage_1_comp_out[67]=i_stage_1_comp_in[32];
assign o_stage_1_comp_out[68]=i_stage_1_comp_in[33];
assign o_stage_1_comp_out[69]=i_stage_1_comp_in[33];
assign o_stage_1_comp_out[70]=i_stage_1_comp_in[33];
assign o_stage_1_comp_out[71]=i_stage_1_comp_in[33];
assign o_stage_1_comp_out[72]=i_stage_1_comp_in[34];
assign o_stage_1_comp_out[73]=i_stage_1_comp_in[34];
assign o_stage_1_comp_out[74]=i_stage_1_comp_in[34];
assign o_stage_1_comp_out[75]=i_stage_1_comp_in[34];
assign o_stage_1_comp_out[76]=i_stage_1_comp_in[35]^i_stage_1_comp_in[36]^i_stage_1_comp_in[37];
assign o_stage_1_comp_out[77]=i_stage_1_comp_in[35]^i_stage_1_comp_in[37];
assign o_stage_1_comp_out[78]=i_stage_1_comp_in[36]^i_stage_1_comp_in[37];
assign o_stage_1_comp_out[79]=i_stage_1_comp_in[37];
assign o_stage_1_comp_out[80]=i_stage_1_comp_in[38];
assign o_stage_1_comp_out[81]=i_stage_1_comp_in[38];
assign o_stage_1_comp_out[82]=i_stage_1_comp_in[38];
assign o_stage_1_comp_out[83]=i_stage_1_comp_in[38];
assign o_stage_1_comp_out[84]=i_stage_1_comp_in[39]^i_stage_1_comp_in[40]^i_stage_1_comp_in[41];
assign o_stage_1_comp_out[85]=i_stage_1_comp_in[39]^i_stage_1_comp_in[41];
assign o_stage_1_comp_out[86]=i_stage_1_comp_in[40]^i_stage_1_comp_in[41];
assign o_stage_1_comp_out[87]=i_stage_1_comp_in[41];
assign o_stage_1_comp_out[88]=i_stage_1_comp_in[42]^i_stage_1_comp_in[43]^i_stage_1_comp_in[44]^i_stage_1_comp_in[45];
assign o_stage_1_comp_out[89]=i_stage_1_comp_in[43]^i_stage_1_comp_in[45];
assign o_stage_1_comp_out[90]=i_stage_1_comp_in[44]^i_stage_1_comp_in[45];
assign o_stage_1_comp_out[91]=i_stage_1_comp_in[45];
assign o_stage_1_comp_out[92]=i_stage_1_comp_in[46]^i_stage_1_comp_in[47]^i_stage_1_comp_in[48]^i_stage_1_comp_in[49];
assign o_stage_1_comp_out[93]=i_stage_1_comp_in[47]^i_stage_1_comp_in[49];
assign o_stage_1_comp_out[94]=i_stage_1_comp_in[48]^i_stage_1_comp_in[49];
assign o_stage_1_comp_out[95]=i_stage_1_comp_in[49];
assign o_stage_1_comp_out[96]=i_stage_1_comp_in[50];
assign o_stage_1_comp_out[97]=i_stage_1_comp_in[50];
assign o_stage_1_comp_out[98]=i_stage_1_comp_in[50];
assign o_stage_1_comp_out[99]=i_stage_1_comp_in[50];
assign o_stage_1_comp_out[100]=i_stage_1_comp_in[51]^i_stage_1_comp_in[52]^i_stage_1_comp_in[53]^i_stage_1_comp_in[54];
assign o_stage_1_comp_out[101]=i_stage_1_comp_in[52]^i_stage_1_comp_in[54];
assign o_stage_1_comp_out[102]=i_stage_1_comp_in[53]^i_stage_1_comp_in[54];
assign o_stage_1_comp_out[103]=i_stage_1_comp_in[54];
assign o_stage_1_comp_out[104]=i_stage_1_comp_in[55]^i_stage_1_comp_in[56]^i_stage_1_comp_in[57]^i_stage_1_comp_in[58];
assign o_stage_1_comp_out[105]=i_stage_1_comp_in[56]^i_stage_1_comp_in[58];
assign o_stage_1_comp_out[106]=i_stage_1_comp_in[57]^i_stage_1_comp_in[58];
assign o_stage_1_comp_out[107]=i_stage_1_comp_in[58];
assign o_stage_1_comp_out[108]=i_stage_1_comp_in[59]^i_stage_1_comp_in[60]^i_stage_1_comp_in[61]^i_stage_1_comp_in[62];
assign o_stage_1_comp_out[109]=i_stage_1_comp_in[60]^i_stage_1_comp_in[62];
assign o_stage_1_comp_out[110]=i_stage_1_comp_in[61]^i_stage_1_comp_in[62];
assign o_stage_1_comp_out[111]=i_stage_1_comp_in[62];
assign o_stage_1_comp_out[112]=i_stage_1_comp_in[63]^i_stage_1_comp_in[64]^i_stage_1_comp_in[65]^i_stage_1_comp_in[66];
assign o_stage_1_comp_out[113]=i_stage_1_comp_in[64]^i_stage_1_comp_in[66];
assign o_stage_1_comp_out[114]=i_stage_1_comp_in[65]^i_stage_1_comp_in[66];
assign o_stage_1_comp_out[115]=i_stage_1_comp_in[66];
assign o_stage_1_comp_out[116]=i_stage_1_comp_in[67]^i_stage_1_comp_in[68]^i_stage_1_comp_in[69]^i_stage_1_comp_in[70];
assign o_stage_1_comp_out[117]=i_stage_1_comp_in[68]^i_stage_1_comp_in[70];
assign o_stage_1_comp_out[118]=i_stage_1_comp_in[69]^i_stage_1_comp_in[70];
assign o_stage_1_comp_out[119]=i_stage_1_comp_in[70];
assign o_stage_1_comp_out[120]=i_stage_1_comp_in[71]^i_stage_1_comp_in[72]^i_stage_1_comp_in[73]^i_stage_1_comp_in[74];
assign o_stage_1_comp_out[121]=i_stage_1_comp_in[72]^i_stage_1_comp_in[74];
assign o_stage_1_comp_out[122]=i_stage_1_comp_in[73]^i_stage_1_comp_in[74];
assign o_stage_1_comp_out[123]=i_stage_1_comp_in[74];
assign o_stage_1_comp_out[124]=i_stage_1_comp_in[75]^i_stage_1_comp_in[76]^i_stage_1_comp_in[77]^i_stage_1_comp_in[78];
assign o_stage_1_comp_out[125]=i_stage_1_comp_in[76]^i_stage_1_comp_in[78];
assign o_stage_1_comp_out[126]=i_stage_1_comp_in[77]^i_stage_1_comp_in[78];
assign o_stage_1_comp_out[127]=i_stage_1_comp_in[78];
assign o_stage_1_comp_out[128]=i_stage_1_comp_in[79];
assign o_stage_1_comp_out[129]=i_stage_1_comp_in[79];
assign o_stage_1_comp_out[130]=i_stage_1_comp_in[79];
assign o_stage_1_comp_out[131]=i_stage_1_comp_in[79];
assign o_stage_1_comp_out[132]=i_stage_1_comp_in[80]^i_stage_1_comp_in[81];
assign o_stage_1_comp_out[133]=i_stage_1_comp_in[81];
assign o_stage_1_comp_out[134]=i_stage_1_comp_in[80]^i_stage_1_comp_in[81];
assign o_stage_1_comp_out[135]=i_stage_1_comp_in[81];
assign o_stage_1_comp_out[136]=i_stage_1_comp_in[82];
assign o_stage_1_comp_out[137]=i_stage_1_comp_in[82];
assign o_stage_1_comp_out[138]=i_stage_1_comp_in[82];
assign o_stage_1_comp_out[139]=i_stage_1_comp_in[82];
assign o_stage_1_comp_out[140]=i_stage_1_comp_in[83]^i_stage_1_comp_in[84]^i_stage_1_comp_in[85];
assign o_stage_1_comp_out[141]=i_stage_1_comp_in[83]^i_stage_1_comp_in[85];
assign o_stage_1_comp_out[142]=i_stage_1_comp_in[84]^i_stage_1_comp_in[85];
assign o_stage_1_comp_out[143]=i_stage_1_comp_in[85];
assign o_stage_1_comp_out[144]=i_stage_1_comp_in[86];
assign o_stage_1_comp_out[145]=i_stage_1_comp_in[86];
assign o_stage_1_comp_out[146]=i_stage_1_comp_in[86];
assign o_stage_1_comp_out[147]=i_stage_1_comp_in[86];
assign o_stage_1_comp_out[148]=i_stage_1_comp_in[87]^i_stage_1_comp_in[88]^i_stage_1_comp_in[89];
assign o_stage_1_comp_out[149]=i_stage_1_comp_in[87]^i_stage_1_comp_in[89];
assign o_stage_1_comp_out[150]=i_stage_1_comp_in[88]^i_stage_1_comp_in[89];
assign o_stage_1_comp_out[151]=i_stage_1_comp_in[89];
assign o_stage_1_comp_out[152]=i_stage_1_comp_in[90]^i_stage_1_comp_in[91]^i_stage_1_comp_in[92];
assign o_stage_1_comp_out[153]=i_stage_1_comp_in[90]^i_stage_1_comp_in[92];
assign o_stage_1_comp_out[154]=i_stage_1_comp_in[91]^i_stage_1_comp_in[92];
assign o_stage_1_comp_out[155]=i_stage_1_comp_in[92];
assign o_stage_1_comp_out[156]=i_stage_1_comp_in[93]^i_stage_1_comp_in[94]^i_stage_1_comp_in[95]^i_stage_1_comp_in[96];
assign o_stage_1_comp_out[157]=i_stage_1_comp_in[94]^i_stage_1_comp_in[96];
assign o_stage_1_comp_out[158]=i_stage_1_comp_in[95]^i_stage_1_comp_in[96];
assign o_stage_1_comp_out[159]=i_stage_1_comp_in[96];
assign o_stage_1_comp_out[160]=i_stage_1_comp_in[97];
assign o_stage_1_comp_out[161]=i_stage_1_comp_in[97];
assign o_stage_1_comp_out[162]=i_stage_1_comp_in[97];
assign o_stage_1_comp_out[163]=i_stage_1_comp_in[97];
assign o_stage_1_comp_out[164]=i_stage_1_comp_in[98];
assign o_stage_1_comp_out[165]=i_stage_1_comp_in[98];
assign o_stage_1_comp_out[166]=i_stage_1_comp_in[98];
assign o_stage_1_comp_out[167]=i_stage_1_comp_in[98];
assign o_stage_1_comp_out[168]=i_stage_1_comp_in[99]^i_stage_1_comp_in[100]^i_stage_1_comp_in[101];
assign o_stage_1_comp_out[169]=i_stage_1_comp_in[99]^i_stage_1_comp_in[101];
assign o_stage_1_comp_out[170]=i_stage_1_comp_in[100]^i_stage_1_comp_in[101];
assign o_stage_1_comp_out[171]=i_stage_1_comp_in[101];
assign o_stage_1_comp_out[172]=i_stage_1_comp_in[102];
assign o_stage_1_comp_out[173]=i_stage_1_comp_in[102];
assign o_stage_1_comp_out[174]=i_stage_1_comp_in[102];
assign o_stage_1_comp_out[175]=i_stage_1_comp_in[102];
assign o_stage_1_comp_out[176]=i_stage_1_comp_in[103];
assign o_stage_1_comp_out[177]=i_stage_1_comp_in[103];
assign o_stage_1_comp_out[178]=i_stage_1_comp_in[103];
assign o_stage_1_comp_out[179]=i_stage_1_comp_in[103];
assign o_stage_1_comp_out[180]=i_stage_1_comp_in[104]^i_stage_1_comp_in[105]^i_stage_1_comp_in[106];
assign o_stage_1_comp_out[181]=i_stage_1_comp_in[104]^i_stage_1_comp_in[106];
assign o_stage_1_comp_out[182]=i_stage_1_comp_in[105]^i_stage_1_comp_in[106];
assign o_stage_1_comp_out[183]=i_stage_1_comp_in[106];
assign o_stage_1_comp_out[184]=i_stage_1_comp_in[107];
assign o_stage_1_comp_out[185]=i_stage_1_comp_in[107];
assign o_stage_1_comp_out[186]=i_stage_1_comp_in[107];
assign o_stage_1_comp_out[187]=i_stage_1_comp_in[107];
assign o_stage_1_comp_out[188]=i_stage_1_comp_in[108]^i_stage_1_comp_in[109]^i_stage_1_comp_in[110]^i_stage_1_comp_in[111];
assign o_stage_1_comp_out[189]=i_stage_1_comp_in[109]^i_stage_1_comp_in[111];
assign o_stage_1_comp_out[190]=i_stage_1_comp_in[110]^i_stage_1_comp_in[111];
assign o_stage_1_comp_out[191]=i_stage_1_comp_in[111];
assign o_stage_1_comp_out[192]=i_stage_1_comp_in[112]^i_stage_1_comp_in[113]^i_stage_1_comp_in[114]^i_stage_1_comp_in[115];
assign o_stage_1_comp_out[193]=i_stage_1_comp_in[113]^i_stage_1_comp_in[115];
assign o_stage_1_comp_out[194]=i_stage_1_comp_in[114]^i_stage_1_comp_in[115];
assign o_stage_1_comp_out[195]=i_stage_1_comp_in[115];
assign o_stage_1_comp_out[196]=i_stage_1_comp_in[116]^i_stage_1_comp_in[117]^i_stage_1_comp_in[118]^i_stage_1_comp_in[119];
assign o_stage_1_comp_out[197]=i_stage_1_comp_in[117]^i_stage_1_comp_in[119];
assign o_stage_1_comp_out[198]=i_stage_1_comp_in[118]^i_stage_1_comp_in[119];
assign o_stage_1_comp_out[199]=i_stage_1_comp_in[119];
assign o_stage_1_comp_out[200]=i_stage_1_comp_in[120];
assign o_stage_1_comp_out[201]=i_stage_1_comp_in[120];
assign o_stage_1_comp_out[202]=i_stage_1_comp_in[120];
assign o_stage_1_comp_out[203]=i_stage_1_comp_in[120];
assign o_stage_1_comp_out[204]=i_stage_1_comp_in[121]^i_stage_1_comp_in[122];
assign o_stage_1_comp_out[205]=i_stage_1_comp_in[122];
assign o_stage_1_comp_out[206]=i_stage_1_comp_in[121]^i_stage_1_comp_in[122];
assign o_stage_1_comp_out[207]=i_stage_1_comp_in[122];
assign o_stage_1_comp_out[208]=i_stage_1_comp_in[123]^i_stage_1_comp_in[124]^i_stage_1_comp_in[125]^i_stage_1_comp_in[126];
assign o_stage_1_comp_out[209]=i_stage_1_comp_in[124]^i_stage_1_comp_in[126];
assign o_stage_1_comp_out[210]=i_stage_1_comp_in[125]^i_stage_1_comp_in[126];
assign o_stage_1_comp_out[211]=i_stage_1_comp_in[126];
assign o_stage_1_comp_out[212]=i_stage_1_comp_in[127]^i_stage_1_comp_in[128]^i_stage_1_comp_in[129];
assign o_stage_1_comp_out[213]=i_stage_1_comp_in[127]^i_stage_1_comp_in[129];
assign o_stage_1_comp_out[214]=i_stage_1_comp_in[128]^i_stage_1_comp_in[129];
assign o_stage_1_comp_out[215]=i_stage_1_comp_in[129];
assign o_stage_1_comp_out[216]=i_stage_1_comp_in[130]^i_stage_1_comp_in[131]^i_stage_1_comp_in[132]^i_stage_1_comp_in[133];
assign o_stage_1_comp_out[217]=i_stage_1_comp_in[131]^i_stage_1_comp_in[133];
assign o_stage_1_comp_out[218]=i_stage_1_comp_in[132]^i_stage_1_comp_in[133];
assign o_stage_1_comp_out[219]=i_stage_1_comp_in[133];
assign o_stage_1_comp_out[220]=i_stage_1_comp_in[134]^i_stage_1_comp_in[135]^i_stage_1_comp_in[136]^i_stage_1_comp_in[137];
assign o_stage_1_comp_out[221]=i_stage_1_comp_in[135]^i_stage_1_comp_in[137];
assign o_stage_1_comp_out[222]=i_stage_1_comp_in[136]^i_stage_1_comp_in[137];
assign o_stage_1_comp_out[223]=i_stage_1_comp_in[137];
assign o_stage_1_comp_out[224]=i_stage_1_comp_in[138]^i_stage_1_comp_in[139]^i_stage_1_comp_in[140]^i_stage_1_comp_in[141];
assign o_stage_1_comp_out[225]=i_stage_1_comp_in[139]^i_stage_1_comp_in[141];
assign o_stage_1_comp_out[226]=i_stage_1_comp_in[140]^i_stage_1_comp_in[141];
assign o_stage_1_comp_out[227]=i_stage_1_comp_in[141];
assign o_stage_1_comp_out[228]=i_stage_1_comp_in[142]^i_stage_1_comp_in[143]^i_stage_1_comp_in[144];
assign o_stage_1_comp_out[229]=i_stage_1_comp_in[142]^i_stage_1_comp_in[144];
assign o_stage_1_comp_out[230]=i_stage_1_comp_in[143]^i_stage_1_comp_in[144];
assign o_stage_1_comp_out[231]=i_stage_1_comp_in[144];
assign o_stage_1_comp_out[232]=i_stage_1_comp_in[145]^i_stage_1_comp_in[146]^i_stage_1_comp_in[147]^i_stage_1_comp_in[148];
assign o_stage_1_comp_out[233]=i_stage_1_comp_in[146]^i_stage_1_comp_in[148];
assign o_stage_1_comp_out[234]=i_stage_1_comp_in[147]^i_stage_1_comp_in[148];
assign o_stage_1_comp_out[235]=i_stage_1_comp_in[148];
assign o_stage_1_comp_out[236]=i_stage_1_comp_in[149]^i_stage_1_comp_in[150]^i_stage_1_comp_in[151]^i_stage_1_comp_in[152];
assign o_stage_1_comp_out[237]=i_stage_1_comp_in[150]^i_stage_1_comp_in[152];
assign o_stage_1_comp_out[238]=i_stage_1_comp_in[151]^i_stage_1_comp_in[152];
assign o_stage_1_comp_out[239]=i_stage_1_comp_in[152];
assign o_stage_1_comp_out[240]=i_stage_1_comp_in[153]^i_stage_1_comp_in[154]^i_stage_1_comp_in[155]^i_stage_1_comp_in[156];
assign o_stage_1_comp_out[241]=i_stage_1_comp_in[154]^i_stage_1_comp_in[156];
assign o_stage_1_comp_out[242]=i_stage_1_comp_in[155]^i_stage_1_comp_in[156];
assign o_stage_1_comp_out[243]=i_stage_1_comp_in[156];
assign o_stage_1_comp_out[244]=i_stage_1_comp_in[157]^i_stage_1_comp_in[158]^i_stage_1_comp_in[159]^i_stage_1_comp_in[160];
assign o_stage_1_comp_out[245]=i_stage_1_comp_in[158]^i_stage_1_comp_in[160];
assign o_stage_1_comp_out[246]=i_stage_1_comp_in[159]^i_stage_1_comp_in[160];
assign o_stage_1_comp_out[247]=i_stage_1_comp_in[160];
assign o_stage_1_comp_out[248]=i_stage_1_comp_in[161]^i_stage_1_comp_in[162]^i_stage_1_comp_in[163]^i_stage_1_comp_in[164];
assign o_stage_1_comp_out[249]=i_stage_1_comp_in[162]^i_stage_1_comp_in[164];
assign o_stage_1_comp_out[250]=i_stage_1_comp_in[163]^i_stage_1_comp_in[164];
assign o_stage_1_comp_out[251]=i_stage_1_comp_in[164];
assign o_stage_1_comp_out[252]=i_stage_1_comp_in[165]^i_stage_1_comp_in[166]^i_stage_1_comp_in[167]^i_stage_1_comp_in[168];
assign o_stage_1_comp_out[253]=i_stage_1_comp_in[166]^i_stage_1_comp_in[168];
assign o_stage_1_comp_out[254]=i_stage_1_comp_in[167]^i_stage_1_comp_in[168];
assign o_stage_1_comp_out[255]=i_stage_1_comp_in[168];
assign o_stage_1_comp_out[256]=i_stage_1_comp_in[169]^i_stage_1_comp_in[170]^i_stage_1_comp_in[171]^i_stage_1_comp_in[172];
assign o_stage_1_comp_out[257]=i_stage_1_comp_in[170]^i_stage_1_comp_in[172];
assign o_stage_1_comp_out[258]=i_stage_1_comp_in[171]^i_stage_1_comp_in[172];
assign o_stage_1_comp_out[259]=i_stage_1_comp_in[172];
assign o_stage_1_comp_out[260]=i_stage_1_comp_in[173];
assign o_stage_1_comp_out[261]=i_stage_1_comp_in[173];
assign o_stage_1_comp_out[262]=i_stage_1_comp_in[173];
assign o_stage_1_comp_out[263]=i_stage_1_comp_in[173];
assign o_stage_1_comp_out[264]=i_stage_1_comp_in[174];
assign o_stage_1_comp_out[265]=i_stage_1_comp_in[174];
assign o_stage_1_comp_out[266]=i_stage_1_comp_in[174];
assign o_stage_1_comp_out[267]=i_stage_1_comp_in[174];
assign o_stage_1_comp_out[268]=i_stage_1_comp_in[175];
assign o_stage_1_comp_out[269]=i_stage_1_comp_in[175];
assign o_stage_1_comp_out[270]=i_stage_1_comp_in[175];
assign o_stage_1_comp_out[271]=i_stage_1_comp_in[175];
assign o_stage_1_comp_out[272]=i_stage_1_comp_in[176]^i_stage_1_comp_in[177]^i_stage_1_comp_in[178]^i_stage_1_comp_in[179];
assign o_stage_1_comp_out[273]=i_stage_1_comp_in[177]^i_stage_1_comp_in[179];
assign o_stage_1_comp_out[274]=i_stage_1_comp_in[178]^i_stage_1_comp_in[179];
assign o_stage_1_comp_out[275]=i_stage_1_comp_in[179];
assign o_stage_1_comp_out[276]=i_stage_1_comp_in[180];
assign o_stage_1_comp_out[277]=i_stage_1_comp_in[180];
assign o_stage_1_comp_out[278]=i_stage_1_comp_in[180];
assign o_stage_1_comp_out[279]=i_stage_1_comp_in[180];
assign o_stage_1_comp_out[280]=i_stage_1_comp_in[181]^i_stage_1_comp_in[182]^i_stage_1_comp_in[183];
assign o_stage_1_comp_out[281]=i_stage_1_comp_in[181]^i_stage_1_comp_in[183];
assign o_stage_1_comp_out[282]=i_stage_1_comp_in[182]^i_stage_1_comp_in[183];
assign o_stage_1_comp_out[283]=i_stage_1_comp_in[183];
assign o_stage_1_comp_out[284]=i_stage_1_comp_in[184]^i_stage_1_comp_in[185]^i_stage_1_comp_in[186]^i_stage_1_comp_in[187];
assign o_stage_1_comp_out[285]=i_stage_1_comp_in[185]^i_stage_1_comp_in[187];
assign o_stage_1_comp_out[286]=i_stage_1_comp_in[186]^i_stage_1_comp_in[187];
assign o_stage_1_comp_out[287]=i_stage_1_comp_in[187];
assign o_stage_1_comp_out[288]=i_stage_1_comp_in[188]^i_stage_1_comp_in[189]^i_stage_1_comp_in[190];
assign o_stage_1_comp_out[289]=i_stage_1_comp_in[188]^i_stage_1_comp_in[190];
assign o_stage_1_comp_out[290]=i_stage_1_comp_in[189]^i_stage_1_comp_in[190];
assign o_stage_1_comp_out[291]=i_stage_1_comp_in[190];
assign o_stage_1_comp_out[292]=i_stage_1_comp_in[191]^i_stage_1_comp_in[192]^i_stage_1_comp_in[193]^i_stage_1_comp_in[194];
assign o_stage_1_comp_out[293]=i_stage_1_comp_in[192]^i_stage_1_comp_in[194];
assign o_stage_1_comp_out[294]=i_stage_1_comp_in[193]^i_stage_1_comp_in[194];
assign o_stage_1_comp_out[295]=i_stage_1_comp_in[194];
assign o_stage_1_comp_out[296]=i_stage_1_comp_in[195]^i_stage_1_comp_in[196]^i_stage_1_comp_in[197]^i_stage_1_comp_in[198];
assign o_stage_1_comp_out[297]=i_stage_1_comp_in[196]^i_stage_1_comp_in[198];
assign o_stage_1_comp_out[298]=i_stage_1_comp_in[197]^i_stage_1_comp_in[198];
assign o_stage_1_comp_out[299]=i_stage_1_comp_in[198];
assign o_stage_1_comp_out[300]=i_stage_1_comp_in[199]^i_stage_1_comp_in[200]^i_stage_1_comp_in[201]^i_stage_1_comp_in[202];
assign o_stage_1_comp_out[301]=i_stage_1_comp_in[200]^i_stage_1_comp_in[202];
assign o_stage_1_comp_out[302]=i_stage_1_comp_in[201]^i_stage_1_comp_in[202];
assign o_stage_1_comp_out[303]=i_stage_1_comp_in[202];
assign o_stage_1_comp_out[304]=i_stage_1_comp_in[203];
assign o_stage_1_comp_out[305]=i_stage_1_comp_in[203];
assign o_stage_1_comp_out[306]=i_stage_1_comp_in[203];
assign o_stage_1_comp_out[307]=i_stage_1_comp_in[203];
assign o_stage_1_comp_out[308]=i_stage_1_comp_in[204]^i_stage_1_comp_in[205]^i_stage_1_comp_in[206];
assign o_stage_1_comp_out[309]=i_stage_1_comp_in[204]^i_stage_1_comp_in[206];
assign o_stage_1_comp_out[310]=i_stage_1_comp_in[205]^i_stage_1_comp_in[206];
assign o_stage_1_comp_out[311]=i_stage_1_comp_in[206];
assign o_stage_1_comp_out[312]=i_stage_1_comp_in[207]^i_stage_1_comp_in[208]^i_stage_1_comp_in[209];
assign o_stage_1_comp_out[313]=i_stage_1_comp_in[207]^i_stage_1_comp_in[209];
assign o_stage_1_comp_out[314]=i_stage_1_comp_in[208]^i_stage_1_comp_in[209];
assign o_stage_1_comp_out[315]=i_stage_1_comp_in[209];
assign o_stage_1_comp_out[316]=i_stage_1_comp_in[210]^i_stage_1_comp_in[211]^i_stage_1_comp_in[212]^i_stage_1_comp_in[213];
assign o_stage_1_comp_out[317]=i_stage_1_comp_in[211]^i_stage_1_comp_in[213];
assign o_stage_1_comp_out[318]=i_stage_1_comp_in[212]^i_stage_1_comp_in[213];
assign o_stage_1_comp_out[319]=i_stage_1_comp_in[213];
assign o_stage_1_comp_out[320]=i_stage_1_comp_in[214]^i_stage_1_comp_in[215]^i_stage_1_comp_in[216];
assign o_stage_1_comp_out[321]=i_stage_1_comp_in[214]^i_stage_1_comp_in[216];
assign o_stage_1_comp_out[322]=i_stage_1_comp_in[215]^i_stage_1_comp_in[216];
assign o_stage_1_comp_out[323]=i_stage_1_comp_in[216];
assign o_stage_1_comp_out[324]=i_stage_1_comp_in[217]^i_stage_1_comp_in[218]^i_stage_1_comp_in[219]^i_stage_1_comp_in[220];
assign o_stage_1_comp_out[325]=i_stage_1_comp_in[218]^i_stage_1_comp_in[220];
assign o_stage_1_comp_out[326]=i_stage_1_comp_in[219]^i_stage_1_comp_in[220];
assign o_stage_1_comp_out[327]=i_stage_1_comp_in[220];
assign o_stage_1_comp_out[328]=i_stage_1_comp_in[221]^i_stage_1_comp_in[222]^i_stage_1_comp_in[223]^i_stage_1_comp_in[224];
assign o_stage_1_comp_out[329]=i_stage_1_comp_in[222]^i_stage_1_comp_in[224];
assign o_stage_1_comp_out[330]=i_stage_1_comp_in[223]^i_stage_1_comp_in[224];
assign o_stage_1_comp_out[331]=i_stage_1_comp_in[224];
assign o_stage_1_comp_out[332]=i_stage_1_comp_in[225]^i_stage_1_comp_in[226]^i_stage_1_comp_in[227]^i_stage_1_comp_in[228];
assign o_stage_1_comp_out[333]=i_stage_1_comp_in[226]^i_stage_1_comp_in[228];
assign o_stage_1_comp_out[334]=i_stage_1_comp_in[227]^i_stage_1_comp_in[228];
assign o_stage_1_comp_out[335]=i_stage_1_comp_in[228];
assign o_stage_1_comp_out[336]=i_stage_1_comp_in[229]^i_stage_1_comp_in[230]^i_stage_1_comp_in[231]^i_stage_1_comp_in[232];
assign o_stage_1_comp_out[337]=i_stage_1_comp_in[230]^i_stage_1_comp_in[232];
assign o_stage_1_comp_out[338]=i_stage_1_comp_in[231]^i_stage_1_comp_in[232];
assign o_stage_1_comp_out[339]=i_stage_1_comp_in[232];
assign o_stage_1_comp_out[340]=i_stage_1_comp_in[233]^i_stage_1_comp_in[234]^i_stage_1_comp_in[235]^i_stage_1_comp_in[236];
assign o_stage_1_comp_out[341]=i_stage_1_comp_in[234]^i_stage_1_comp_in[236];
assign o_stage_1_comp_out[342]=i_stage_1_comp_in[235]^i_stage_1_comp_in[236];
assign o_stage_1_comp_out[343]=i_stage_1_comp_in[236];
assign o_stage_1_comp_out[344]=i_stage_1_comp_in[237]^i_stage_1_comp_in[238]^i_stage_1_comp_in[239]^i_stage_1_comp_in[240];
assign o_stage_1_comp_out[345]=i_stage_1_comp_in[238]^i_stage_1_comp_in[240];
assign o_stage_1_comp_out[346]=i_stage_1_comp_in[239]^i_stage_1_comp_in[240];
assign o_stage_1_comp_out[347]=i_stage_1_comp_in[240];
assign o_stage_1_comp_out[348]=i_stage_1_comp_in[241]^i_stage_1_comp_in[242]^i_stage_1_comp_in[243]^i_stage_1_comp_in[244];
assign o_stage_1_comp_out[349]=i_stage_1_comp_in[242]^i_stage_1_comp_in[244];
assign o_stage_1_comp_out[350]=i_stage_1_comp_in[243]^i_stage_1_comp_in[244];
assign o_stage_1_comp_out[351]=i_stage_1_comp_in[244];
assign o_stage_1_comp_out[352]=i_stage_1_comp_in[245]^i_stage_1_comp_in[246]^i_stage_1_comp_in[247]^i_stage_1_comp_in[248];
assign o_stage_1_comp_out[353]=i_stage_1_comp_in[246]^i_stage_1_comp_in[248];
assign o_stage_1_comp_out[354]=i_stage_1_comp_in[247]^i_stage_1_comp_in[248];
assign o_stage_1_comp_out[355]=i_stage_1_comp_in[248];
assign o_stage_1_comp_out[356]=i_stage_1_comp_in[249]^i_stage_1_comp_in[250]^i_stage_1_comp_in[251]^i_stage_1_comp_in[252];
assign o_stage_1_comp_out[357]=i_stage_1_comp_in[250]^i_stage_1_comp_in[252];
assign o_stage_1_comp_out[358]=i_stage_1_comp_in[251]^i_stage_1_comp_in[252];
assign o_stage_1_comp_out[359]=i_stage_1_comp_in[252];
assign o_stage_1_comp_out[360]=i_stage_1_comp_in[253]^i_stage_1_comp_in[254]^i_stage_1_comp_in[255]^i_stage_1_comp_in[256];
assign o_stage_1_comp_out[361]=i_stage_1_comp_in[254]^i_stage_1_comp_in[256];
assign o_stage_1_comp_out[362]=i_stage_1_comp_in[255]^i_stage_1_comp_in[256];
assign o_stage_1_comp_out[363]=i_stage_1_comp_in[256];
assign o_stage_1_comp_out[364]=i_stage_1_comp_in[257]^i_stage_1_comp_in[258]^i_stage_1_comp_in[259]^i_stage_1_comp_in[260];
assign o_stage_1_comp_out[365]=i_stage_1_comp_in[258]^i_stage_1_comp_in[260];
assign o_stage_1_comp_out[366]=i_stage_1_comp_in[259]^i_stage_1_comp_in[260];
assign o_stage_1_comp_out[367]=i_stage_1_comp_in[260];
assign o_stage_1_comp_out[368]=i_stage_1_comp_in[261];
assign o_stage_1_comp_out[369]=i_stage_1_comp_in[261];
assign o_stage_1_comp_out[370]=i_stage_1_comp_in[261];
assign o_stage_1_comp_out[371]=i_stage_1_comp_in[261];
assign o_stage_1_comp_out[372]=i_stage_1_comp_in[262]^i_stage_1_comp_in[263]^i_stage_1_comp_in[264];
assign o_stage_1_comp_out[373]=i_stage_1_comp_in[262]^i_stage_1_comp_in[264];
assign o_stage_1_comp_out[374]=i_stage_1_comp_in[263]^i_stage_1_comp_in[264];
assign o_stage_1_comp_out[375]=i_stage_1_comp_in[264];
assign o_stage_1_comp_out[376]=i_stage_1_comp_in[265]^i_stage_1_comp_in[266]^i_stage_1_comp_in[267];
assign o_stage_1_comp_out[377]=i_stage_1_comp_in[265]^i_stage_1_comp_in[267];
assign o_stage_1_comp_out[378]=i_stage_1_comp_in[266]^i_stage_1_comp_in[267];
assign o_stage_1_comp_out[379]=i_stage_1_comp_in[267];
assign o_stage_1_comp_out[380]=i_stage_1_comp_in[268]^i_stage_1_comp_in[269]^i_stage_1_comp_in[270]^i_stage_1_comp_in[271];
assign o_stage_1_comp_out[381]=i_stage_1_comp_in[269]^i_stage_1_comp_in[271];
assign o_stage_1_comp_out[382]=i_stage_1_comp_in[270]^i_stage_1_comp_in[271];
assign o_stage_1_comp_out[383]=i_stage_1_comp_in[271];
assign o_stage_1_comp_out[384]=i_stage_1_comp_in[272]^i_stage_1_comp_in[273]^i_stage_1_comp_in[274]^i_stage_1_comp_in[275];
assign o_stage_1_comp_out[385]=i_stage_1_comp_in[273]^i_stage_1_comp_in[275];
assign o_stage_1_comp_out[386]=i_stage_1_comp_in[274]^i_stage_1_comp_in[275];
assign o_stage_1_comp_out[387]=i_stage_1_comp_in[275];
assign o_stage_1_comp_out[388]=i_stage_1_comp_in[276]^i_stage_1_comp_in[277]^i_stage_1_comp_in[278]^i_stage_1_comp_in[279];
assign o_stage_1_comp_out[389]=i_stage_1_comp_in[277]^i_stage_1_comp_in[279];
assign o_stage_1_comp_out[390]=i_stage_1_comp_in[278]^i_stage_1_comp_in[279];
assign o_stage_1_comp_out[391]=i_stage_1_comp_in[279];
assign o_stage_1_comp_out[392]=i_stage_1_comp_in[280]^i_stage_1_comp_in[281]^i_stage_1_comp_in[282]^i_stage_1_comp_in[283];
assign o_stage_1_comp_out[393]=i_stage_1_comp_in[281]^i_stage_1_comp_in[283];
assign o_stage_1_comp_out[394]=i_stage_1_comp_in[282]^i_stage_1_comp_in[283];
assign o_stage_1_comp_out[395]=i_stage_1_comp_in[283];
assign o_stage_1_comp_out[396]=i_stage_1_comp_in[284]^i_stage_1_comp_in[285]^i_stage_1_comp_in[286]^i_stage_1_comp_in[287];
assign o_stage_1_comp_out[397]=i_stage_1_comp_in[285]^i_stage_1_comp_in[287];
assign o_stage_1_comp_out[398]=i_stage_1_comp_in[286]^i_stage_1_comp_in[287];
assign o_stage_1_comp_out[399]=i_stage_1_comp_in[287];
assign o_stage_1_comp_out[400]=i_stage_1_comp_in[288]^i_stage_1_comp_in[289]^i_stage_1_comp_in[290]^i_stage_1_comp_in[291];
assign o_stage_1_comp_out[401]=i_stage_1_comp_in[289]^i_stage_1_comp_in[291];
assign o_stage_1_comp_out[402]=i_stage_1_comp_in[290]^i_stage_1_comp_in[291];
assign o_stage_1_comp_out[403]=i_stage_1_comp_in[291];
assign o_stage_1_comp_out[404]=i_stage_1_comp_in[292]^i_stage_1_comp_in[293]^i_stage_1_comp_in[294]^i_stage_1_comp_in[295];
assign o_stage_1_comp_out[405]=i_stage_1_comp_in[293]^i_stage_1_comp_in[295];
assign o_stage_1_comp_out[406]=i_stage_1_comp_in[294]^i_stage_1_comp_in[295];
assign o_stage_1_comp_out[407]=i_stage_1_comp_in[295];
assign o_stage_1_comp_out[408]=i_stage_1_comp_in[296]^i_stage_1_comp_in[297]^i_stage_1_comp_in[298]^i_stage_1_comp_in[299];
assign o_stage_1_comp_out[409]=i_stage_1_comp_in[297]^i_stage_1_comp_in[299];
assign o_stage_1_comp_out[410]=i_stage_1_comp_in[298]^i_stage_1_comp_in[299];
assign o_stage_1_comp_out[411]=i_stage_1_comp_in[299];
assign o_stage_1_comp_out[412]=i_stage_1_comp_in[300]^i_stage_1_comp_in[301]^i_stage_1_comp_in[302]^i_stage_1_comp_in[303];
assign o_stage_1_comp_out[413]=i_stage_1_comp_in[301]^i_stage_1_comp_in[303];
assign o_stage_1_comp_out[414]=i_stage_1_comp_in[302]^i_stage_1_comp_in[303];
assign o_stage_1_comp_out[415]=i_stage_1_comp_in[303];
assign o_stage_1_comp_out[416]=i_stage_1_comp_in[304]^i_stage_1_comp_in[305]^i_stage_1_comp_in[306]^i_stage_1_comp_in[307];
assign o_stage_1_comp_out[417]=i_stage_1_comp_in[305]^i_stage_1_comp_in[307];
assign o_stage_1_comp_out[418]=i_stage_1_comp_in[306]^i_stage_1_comp_in[307];
assign o_stage_1_comp_out[419]=i_stage_1_comp_in[307];
assign o_stage_1_comp_out[420]=i_stage_1_comp_in[308]^i_stage_1_comp_in[309]^i_stage_1_comp_in[310]^i_stage_1_comp_in[311];
assign o_stage_1_comp_out[421]=i_stage_1_comp_in[309]^i_stage_1_comp_in[311];
assign o_stage_1_comp_out[422]=i_stage_1_comp_in[310]^i_stage_1_comp_in[311];
assign o_stage_1_comp_out[423]=i_stage_1_comp_in[311];
assign o_stage_1_comp_out[424]=i_stage_1_comp_in[312]^i_stage_1_comp_in[313]^i_stage_1_comp_in[314]^i_stage_1_comp_in[315];
assign o_stage_1_comp_out[425]=i_stage_1_comp_in[313]^i_stage_1_comp_in[315];
assign o_stage_1_comp_out[426]=i_stage_1_comp_in[314]^i_stage_1_comp_in[315];
assign o_stage_1_comp_out[427]=i_stage_1_comp_in[315];
assign o_stage_1_comp_out[428]=i_stage_1_comp_in[316]^i_stage_1_comp_in[317]^i_stage_1_comp_in[318]^i_stage_1_comp_in[319];
assign o_stage_1_comp_out[429]=i_stage_1_comp_in[317]^i_stage_1_comp_in[319];
assign o_stage_1_comp_out[430]=i_stage_1_comp_in[318]^i_stage_1_comp_in[319];
assign o_stage_1_comp_out[431]=i_stage_1_comp_in[319];
assign o_stage_1_comp_out[432]=i_stage_1_comp_in[320]^i_stage_1_comp_in[321]^i_stage_1_comp_in[322]^i_stage_1_comp_in[323];
assign o_stage_1_comp_out[433]=i_stage_1_comp_in[321]^i_stage_1_comp_in[323];
assign o_stage_1_comp_out[434]=i_stage_1_comp_in[322]^i_stage_1_comp_in[323];
assign o_stage_1_comp_out[435]=i_stage_1_comp_in[323];
assign o_stage_1_comp_out[436]=i_stage_1_comp_in[324]^i_stage_1_comp_in[325]^i_stage_1_comp_in[326]^i_stage_1_comp_in[327];
assign o_stage_1_comp_out[437]=i_stage_1_comp_in[325]^i_stage_1_comp_in[327];
assign o_stage_1_comp_out[438]=i_stage_1_comp_in[326]^i_stage_1_comp_in[327];
assign o_stage_1_comp_out[439]=i_stage_1_comp_in[327];
assign o_stage_1_comp_out[440]=i_stage_1_comp_in[328]^i_stage_1_comp_in[329]^i_stage_1_comp_in[330]^i_stage_1_comp_in[331];
assign o_stage_1_comp_out[441]=i_stage_1_comp_in[329]^i_stage_1_comp_in[331];
assign o_stage_1_comp_out[442]=i_stage_1_comp_in[330]^i_stage_1_comp_in[331];
assign o_stage_1_comp_out[443]=i_stage_1_comp_in[331];
assign o_stage_1_comp_out[444]=i_stage_1_comp_in[332]^i_stage_1_comp_in[333]^i_stage_1_comp_in[334]^i_stage_1_comp_in[335];
assign o_stage_1_comp_out[445]=i_stage_1_comp_in[333]^i_stage_1_comp_in[335];
assign o_stage_1_comp_out[446]=i_stage_1_comp_in[334]^i_stage_1_comp_in[335];
assign o_stage_1_comp_out[447]=i_stage_1_comp_in[335];
assign o_stage_1_comp_out[448]=i_stage_1_comp_in[336]^i_stage_1_comp_in[337]^i_stage_1_comp_in[338]^i_stage_1_comp_in[339];
assign o_stage_1_comp_out[449]=i_stage_1_comp_in[337]^i_stage_1_comp_in[339];
assign o_stage_1_comp_out[450]=i_stage_1_comp_in[338]^i_stage_1_comp_in[339];
assign o_stage_1_comp_out[451]=i_stage_1_comp_in[339];
assign o_stage_1_comp_out[452]=i_stage_1_comp_in[340]^i_stage_1_comp_in[341]^i_stage_1_comp_in[342]^i_stage_1_comp_in[343];
assign o_stage_1_comp_out[453]=i_stage_1_comp_in[341]^i_stage_1_comp_in[343];
assign o_stage_1_comp_out[454]=i_stage_1_comp_in[342]^i_stage_1_comp_in[343];
assign o_stage_1_comp_out[455]=i_stage_1_comp_in[343];
assign o_stage_1_comp_out[456]=i_stage_1_comp_in[344]^i_stage_1_comp_in[345]^i_stage_1_comp_in[346]^i_stage_1_comp_in[347];
assign o_stage_1_comp_out[457]=i_stage_1_comp_in[345]^i_stage_1_comp_in[347];
assign o_stage_1_comp_out[458]=i_stage_1_comp_in[346]^i_stage_1_comp_in[347];
assign o_stage_1_comp_out[459]=i_stage_1_comp_in[347];
assign o_stage_1_comp_out[460]=i_stage_1_comp_in[348]^i_stage_1_comp_in[349]^i_stage_1_comp_in[350]^i_stage_1_comp_in[351];
assign o_stage_1_comp_out[461]=i_stage_1_comp_in[349]^i_stage_1_comp_in[351];
assign o_stage_1_comp_out[462]=i_stage_1_comp_in[350]^i_stage_1_comp_in[351];
assign o_stage_1_comp_out[463]=i_stage_1_comp_in[351];
assign o_stage_1_comp_out[464]=i_stage_1_comp_in[352]^i_stage_1_comp_in[353]^i_stage_1_comp_in[354]^i_stage_1_comp_in[355];
assign o_stage_1_comp_out[465]=i_stage_1_comp_in[353]^i_stage_1_comp_in[355];
assign o_stage_1_comp_out[466]=i_stage_1_comp_in[354]^i_stage_1_comp_in[355];
assign o_stage_1_comp_out[467]=i_stage_1_comp_in[355];
assign o_stage_1_comp_out[468]=i_stage_1_comp_in[356]^i_stage_1_comp_in[357]^i_stage_1_comp_in[358]^i_stage_1_comp_in[359];
assign o_stage_1_comp_out[469]=i_stage_1_comp_in[357]^i_stage_1_comp_in[359];
assign o_stage_1_comp_out[470]=i_stage_1_comp_in[358]^i_stage_1_comp_in[359];
assign o_stage_1_comp_out[471]=i_stage_1_comp_in[359];
assign o_stage_1_comp_out[472]=i_stage_1_comp_in[360]^i_stage_1_comp_in[361]^i_stage_1_comp_in[362]^i_stage_1_comp_in[363];
assign o_stage_1_comp_out[473]=i_stage_1_comp_in[361]^i_stage_1_comp_in[363];
assign o_stage_1_comp_out[474]=i_stage_1_comp_in[362]^i_stage_1_comp_in[363];
assign o_stage_1_comp_out[475]=i_stage_1_comp_in[363];
assign o_stage_1_comp_out[476]=i_stage_1_comp_in[364]^i_stage_1_comp_in[365]^i_stage_1_comp_in[366]^i_stage_1_comp_in[367];
assign o_stage_1_comp_out[477]=i_stage_1_comp_in[365]^i_stage_1_comp_in[367];
assign o_stage_1_comp_out[478]=i_stage_1_comp_in[366]^i_stage_1_comp_in[367];
assign o_stage_1_comp_out[479]=i_stage_1_comp_in[367];
assign o_stage_1_comp_out[480]=i_stage_1_comp_in[368]^i_stage_1_comp_in[369]^i_stage_1_comp_in[370]^i_stage_1_comp_in[371];
assign o_stage_1_comp_out[481]=i_stage_1_comp_in[369]^i_stage_1_comp_in[371];
assign o_stage_1_comp_out[482]=i_stage_1_comp_in[370]^i_stage_1_comp_in[371];
assign o_stage_1_comp_out[483]=i_stage_1_comp_in[371];
assign o_stage_1_comp_out[484]=i_stage_1_comp_in[372]^i_stage_1_comp_in[373]^i_stage_1_comp_in[374]^i_stage_1_comp_in[375];
assign o_stage_1_comp_out[485]=i_stage_1_comp_in[373]^i_stage_1_comp_in[375];
assign o_stage_1_comp_out[486]=i_stage_1_comp_in[374]^i_stage_1_comp_in[375];
assign o_stage_1_comp_out[487]=i_stage_1_comp_in[375];
assign o_stage_1_comp_out[488]=i_stage_1_comp_in[376]^i_stage_1_comp_in[377]^i_stage_1_comp_in[378]^i_stage_1_comp_in[379];
assign o_stage_1_comp_out[489]=i_stage_1_comp_in[377]^i_stage_1_comp_in[379];
assign o_stage_1_comp_out[490]=i_stage_1_comp_in[378]^i_stage_1_comp_in[379];
assign o_stage_1_comp_out[491]=i_stage_1_comp_in[379];
assign o_stage_1_comp_out[492]=i_stage_1_comp_in[380]^i_stage_1_comp_in[381]^i_stage_1_comp_in[382]^i_stage_1_comp_in[383];
assign o_stage_1_comp_out[493]=i_stage_1_comp_in[381]^i_stage_1_comp_in[383];
assign o_stage_1_comp_out[494]=i_stage_1_comp_in[382]^i_stage_1_comp_in[383];
assign o_stage_1_comp_out[495]=i_stage_1_comp_in[383];


endmodule

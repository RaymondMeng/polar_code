`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/04/05 16:57:45
// Design Name: 
// Module Name: stage_6_xor_unit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`include "defines.v"

module stage_6_xor_unit(
    input [`STAGE6_INPUT_WIDTH-1 : 0] i_stage_6_comp_in,  //compute input
    output [`STAGE6_OUTPUT_WIDTH-1 : 0] o_stage_6_comp_out //compute output
    );

assign o_stage_6_comp_out[0]=i_stage_6_comp_in[0]^i_stage_6_comp_in[512];
assign o_stage_6_comp_out[1]=i_stage_6_comp_in[1]^i_stage_6_comp_in[513];
assign o_stage_6_comp_out[2]=i_stage_6_comp_in[2]^i_stage_6_comp_in[514];
assign o_stage_6_comp_out[3]=i_stage_6_comp_in[3]^i_stage_6_comp_in[515];
assign o_stage_6_comp_out[4]=i_stage_6_comp_in[4]^i_stage_6_comp_in[516];
assign o_stage_6_comp_out[5]=i_stage_6_comp_in[5]^i_stage_6_comp_in[517];
assign o_stage_6_comp_out[6]=i_stage_6_comp_in[6]^i_stage_6_comp_in[518];
assign o_stage_6_comp_out[7]=i_stage_6_comp_in[7]^i_stage_6_comp_in[519];
assign o_stage_6_comp_out[8]=i_stage_6_comp_in[8]^i_stage_6_comp_in[520];
assign o_stage_6_comp_out[9]=i_stage_6_comp_in[9]^i_stage_6_comp_in[521];
assign o_stage_6_comp_out[10]=i_stage_6_comp_in[10]^i_stage_6_comp_in[522];
assign o_stage_6_comp_out[11]=i_stage_6_comp_in[11]^i_stage_6_comp_in[523];
assign o_stage_6_comp_out[12]=i_stage_6_comp_in[12]^i_stage_6_comp_in[524];
assign o_stage_6_comp_out[13]=i_stage_6_comp_in[13]^i_stage_6_comp_in[525];
assign o_stage_6_comp_out[14]=i_stage_6_comp_in[14]^i_stage_6_comp_in[526];
assign o_stage_6_comp_out[15]=i_stage_6_comp_in[15]^i_stage_6_comp_in[527];
assign o_stage_6_comp_out[16]=i_stage_6_comp_in[16]^i_stage_6_comp_in[528];
assign o_stage_6_comp_out[17]=i_stage_6_comp_in[17]^i_stage_6_comp_in[529];
assign o_stage_6_comp_out[18]=i_stage_6_comp_in[18]^i_stage_6_comp_in[530];
assign o_stage_6_comp_out[19]=i_stage_6_comp_in[19]^i_stage_6_comp_in[531];
assign o_stage_6_comp_out[20]=i_stage_6_comp_in[20]^i_stage_6_comp_in[532];
assign o_stage_6_comp_out[21]=i_stage_6_comp_in[21]^i_stage_6_comp_in[533];
assign o_stage_6_comp_out[22]=i_stage_6_comp_in[22]^i_stage_6_comp_in[534];
assign o_stage_6_comp_out[23]=i_stage_6_comp_in[23]^i_stage_6_comp_in[535];
assign o_stage_6_comp_out[24]=i_stage_6_comp_in[24]^i_stage_6_comp_in[536];
assign o_stage_6_comp_out[25]=i_stage_6_comp_in[25]^i_stage_6_comp_in[537];
assign o_stage_6_comp_out[26]=i_stage_6_comp_in[26]^i_stage_6_comp_in[538];
assign o_stage_6_comp_out[27]=i_stage_6_comp_in[27]^i_stage_6_comp_in[539];
assign o_stage_6_comp_out[28]=i_stage_6_comp_in[28]^i_stage_6_comp_in[540];
assign o_stage_6_comp_out[29]=i_stage_6_comp_in[29]^i_stage_6_comp_in[541];
assign o_stage_6_comp_out[30]=i_stage_6_comp_in[30]^i_stage_6_comp_in[542];
assign o_stage_6_comp_out[31]=i_stage_6_comp_in[31]^i_stage_6_comp_in[543];
assign o_stage_6_comp_out[32]=i_stage_6_comp_in[32]^i_stage_6_comp_in[544];
assign o_stage_6_comp_out[33]=i_stage_6_comp_in[33]^i_stage_6_comp_in[545];
assign o_stage_6_comp_out[34]=i_stage_6_comp_in[34]^i_stage_6_comp_in[546];
assign o_stage_6_comp_out[35]=i_stage_6_comp_in[35]^i_stage_6_comp_in[547];
assign o_stage_6_comp_out[36]=i_stage_6_comp_in[36]^i_stage_6_comp_in[548];
assign o_stage_6_comp_out[37]=i_stage_6_comp_in[37]^i_stage_6_comp_in[549];
assign o_stage_6_comp_out[38]=i_stage_6_comp_in[38]^i_stage_6_comp_in[550];
assign o_stage_6_comp_out[39]=i_stage_6_comp_in[39]^i_stage_6_comp_in[551];
assign o_stage_6_comp_out[40]=i_stage_6_comp_in[40]^i_stage_6_comp_in[552];
assign o_stage_6_comp_out[41]=i_stage_6_comp_in[41]^i_stage_6_comp_in[553];
assign o_stage_6_comp_out[42]=i_stage_6_comp_in[42]^i_stage_6_comp_in[554];
assign o_stage_6_comp_out[43]=i_stage_6_comp_in[43]^i_stage_6_comp_in[555];
assign o_stage_6_comp_out[44]=i_stage_6_comp_in[44]^i_stage_6_comp_in[556];
assign o_stage_6_comp_out[45]=i_stage_6_comp_in[45]^i_stage_6_comp_in[557];
assign o_stage_6_comp_out[46]=i_stage_6_comp_in[46]^i_stage_6_comp_in[558];
assign o_stage_6_comp_out[47]=i_stage_6_comp_in[47]^i_stage_6_comp_in[559];
assign o_stage_6_comp_out[48]=i_stage_6_comp_in[48]^i_stage_6_comp_in[560];
assign o_stage_6_comp_out[49]=i_stage_6_comp_in[49]^i_stage_6_comp_in[561];
assign o_stage_6_comp_out[50]=i_stage_6_comp_in[50]^i_stage_6_comp_in[562];
assign o_stage_6_comp_out[51]=i_stage_6_comp_in[51]^i_stage_6_comp_in[563];
assign o_stage_6_comp_out[52]=i_stage_6_comp_in[52]^i_stage_6_comp_in[564];
assign o_stage_6_comp_out[53]=i_stage_6_comp_in[53]^i_stage_6_comp_in[565];
assign o_stage_6_comp_out[54]=i_stage_6_comp_in[54]^i_stage_6_comp_in[566];
assign o_stage_6_comp_out[55]=i_stage_6_comp_in[55]^i_stage_6_comp_in[567];
assign o_stage_6_comp_out[56]=i_stage_6_comp_in[56]^i_stage_6_comp_in[568];
assign o_stage_6_comp_out[57]=i_stage_6_comp_in[57]^i_stage_6_comp_in[569];
assign o_stage_6_comp_out[58]=i_stage_6_comp_in[58]^i_stage_6_comp_in[570];
assign o_stage_6_comp_out[59]=i_stage_6_comp_in[59]^i_stage_6_comp_in[571];
assign o_stage_6_comp_out[60]=i_stage_6_comp_in[60]^i_stage_6_comp_in[572];
assign o_stage_6_comp_out[61]=i_stage_6_comp_in[61]^i_stage_6_comp_in[573];
assign o_stage_6_comp_out[62]=i_stage_6_comp_in[62]^i_stage_6_comp_in[574];
assign o_stage_6_comp_out[63]=i_stage_6_comp_in[63]^i_stage_6_comp_in[575];
assign o_stage_6_comp_out[64]=i_stage_6_comp_in[64]^i_stage_6_comp_in[576];
assign o_stage_6_comp_out[65]=i_stage_6_comp_in[65]^i_stage_6_comp_in[577];
assign o_stage_6_comp_out[66]=i_stage_6_comp_in[66]^i_stage_6_comp_in[578];
assign o_stage_6_comp_out[67]=i_stage_6_comp_in[67]^i_stage_6_comp_in[579];
assign o_stage_6_comp_out[68]=i_stage_6_comp_in[68]^i_stage_6_comp_in[580];
assign o_stage_6_comp_out[69]=i_stage_6_comp_in[69]^i_stage_6_comp_in[581];
assign o_stage_6_comp_out[70]=i_stage_6_comp_in[70]^i_stage_6_comp_in[582];
assign o_stage_6_comp_out[71]=i_stage_6_comp_in[71]^i_stage_6_comp_in[583];
assign o_stage_6_comp_out[72]=i_stage_6_comp_in[72]^i_stage_6_comp_in[584];
assign o_stage_6_comp_out[73]=i_stage_6_comp_in[73]^i_stage_6_comp_in[585];
assign o_stage_6_comp_out[74]=i_stage_6_comp_in[74]^i_stage_6_comp_in[586];
assign o_stage_6_comp_out[75]=i_stage_6_comp_in[75]^i_stage_6_comp_in[587];
assign o_stage_6_comp_out[76]=i_stage_6_comp_in[76]^i_stage_6_comp_in[588];
assign o_stage_6_comp_out[77]=i_stage_6_comp_in[77]^i_stage_6_comp_in[589];
assign o_stage_6_comp_out[78]=i_stage_6_comp_in[78]^i_stage_6_comp_in[590];
assign o_stage_6_comp_out[79]=i_stage_6_comp_in[79]^i_stage_6_comp_in[591];
assign o_stage_6_comp_out[80]=i_stage_6_comp_in[80]^i_stage_6_comp_in[592];
assign o_stage_6_comp_out[81]=i_stage_6_comp_in[81]^i_stage_6_comp_in[593];
assign o_stage_6_comp_out[82]=i_stage_6_comp_in[82]^i_stage_6_comp_in[594];
assign o_stage_6_comp_out[83]=i_stage_6_comp_in[83]^i_stage_6_comp_in[595];
assign o_stage_6_comp_out[84]=i_stage_6_comp_in[84]^i_stage_6_comp_in[596];
assign o_stage_6_comp_out[85]=i_stage_6_comp_in[85]^i_stage_6_comp_in[597];
assign o_stage_6_comp_out[86]=i_stage_6_comp_in[86]^i_stage_6_comp_in[598];
assign o_stage_6_comp_out[87]=i_stage_6_comp_in[87]^i_stage_6_comp_in[599];
assign o_stage_6_comp_out[88]=i_stage_6_comp_in[88]^i_stage_6_comp_in[600];
assign o_stage_6_comp_out[89]=i_stage_6_comp_in[89]^i_stage_6_comp_in[601];
assign o_stage_6_comp_out[90]=i_stage_6_comp_in[90]^i_stage_6_comp_in[602];
assign o_stage_6_comp_out[91]=i_stage_6_comp_in[91]^i_stage_6_comp_in[603];
assign o_stage_6_comp_out[92]=i_stage_6_comp_in[92]^i_stage_6_comp_in[604];
assign o_stage_6_comp_out[93]=i_stage_6_comp_in[93]^i_stage_6_comp_in[605];
assign o_stage_6_comp_out[94]=i_stage_6_comp_in[94]^i_stage_6_comp_in[606];
assign o_stage_6_comp_out[95]=i_stage_6_comp_in[95]^i_stage_6_comp_in[607];
assign o_stage_6_comp_out[96]=i_stage_6_comp_in[96]^i_stage_6_comp_in[608];
assign o_stage_6_comp_out[97]=i_stage_6_comp_in[97]^i_stage_6_comp_in[609];
assign o_stage_6_comp_out[98]=i_stage_6_comp_in[98]^i_stage_6_comp_in[610];
assign o_stage_6_comp_out[99]=i_stage_6_comp_in[99]^i_stage_6_comp_in[611];
assign o_stage_6_comp_out[100]=i_stage_6_comp_in[100]^i_stage_6_comp_in[612];
assign o_stage_6_comp_out[101]=i_stage_6_comp_in[101]^i_stage_6_comp_in[613];
assign o_stage_6_comp_out[102]=i_stage_6_comp_in[102]^i_stage_6_comp_in[614];
assign o_stage_6_comp_out[103]=i_stage_6_comp_in[103]^i_stage_6_comp_in[615];
assign o_stage_6_comp_out[104]=i_stage_6_comp_in[104]^i_stage_6_comp_in[616];
assign o_stage_6_comp_out[105]=i_stage_6_comp_in[105]^i_stage_6_comp_in[617];
assign o_stage_6_comp_out[106]=i_stage_6_comp_in[106]^i_stage_6_comp_in[618];
assign o_stage_6_comp_out[107]=i_stage_6_comp_in[107]^i_stage_6_comp_in[619];
assign o_stage_6_comp_out[108]=i_stage_6_comp_in[108]^i_stage_6_comp_in[620];
assign o_stage_6_comp_out[109]=i_stage_6_comp_in[109]^i_stage_6_comp_in[621];
assign o_stage_6_comp_out[110]=i_stage_6_comp_in[110]^i_stage_6_comp_in[622];
assign o_stage_6_comp_out[111]=i_stage_6_comp_in[111]^i_stage_6_comp_in[623];
assign o_stage_6_comp_out[112]=i_stage_6_comp_in[112]^i_stage_6_comp_in[624];
assign o_stage_6_comp_out[113]=i_stage_6_comp_in[113]^i_stage_6_comp_in[625];
assign o_stage_6_comp_out[114]=i_stage_6_comp_in[114]^i_stage_6_comp_in[626];
assign o_stage_6_comp_out[115]=i_stage_6_comp_in[115]^i_stage_6_comp_in[627];
assign o_stage_6_comp_out[116]=i_stage_6_comp_in[116]^i_stage_6_comp_in[628];
assign o_stage_6_comp_out[117]=i_stage_6_comp_in[117]^i_stage_6_comp_in[629];
assign o_stage_6_comp_out[118]=i_stage_6_comp_in[118]^i_stage_6_comp_in[630];
assign o_stage_6_comp_out[119]=i_stage_6_comp_in[119]^i_stage_6_comp_in[631];
assign o_stage_6_comp_out[120]=i_stage_6_comp_in[120]^i_stage_6_comp_in[632];
assign o_stage_6_comp_out[121]=i_stage_6_comp_in[121]^i_stage_6_comp_in[633];
assign o_stage_6_comp_out[122]=i_stage_6_comp_in[122]^i_stage_6_comp_in[634];
assign o_stage_6_comp_out[123]=i_stage_6_comp_in[123]^i_stage_6_comp_in[635];
assign o_stage_6_comp_out[124]=i_stage_6_comp_in[124]^i_stage_6_comp_in[636];
assign o_stage_6_comp_out[125]=i_stage_6_comp_in[125]^i_stage_6_comp_in[637];
assign o_stage_6_comp_out[126]=i_stage_6_comp_in[126]^i_stage_6_comp_in[638];
assign o_stage_6_comp_out[127]=i_stage_6_comp_in[127]^i_stage_6_comp_in[639];
assign o_stage_6_comp_out[128]=i_stage_6_comp_in[128]^i_stage_6_comp_in[640];
assign o_stage_6_comp_out[129]=i_stage_6_comp_in[129]^i_stage_6_comp_in[641];
assign o_stage_6_comp_out[130]=i_stage_6_comp_in[130]^i_stage_6_comp_in[642];
assign o_stage_6_comp_out[131]=i_stage_6_comp_in[131]^i_stage_6_comp_in[643];
assign o_stage_6_comp_out[132]=i_stage_6_comp_in[132]^i_stage_6_comp_in[644];
assign o_stage_6_comp_out[133]=i_stage_6_comp_in[133]^i_stage_6_comp_in[645];
assign o_stage_6_comp_out[134]=i_stage_6_comp_in[134]^i_stage_6_comp_in[646];
assign o_stage_6_comp_out[135]=i_stage_6_comp_in[135]^i_stage_6_comp_in[647];
assign o_stage_6_comp_out[136]=i_stage_6_comp_in[136]^i_stage_6_comp_in[648];
assign o_stage_6_comp_out[137]=i_stage_6_comp_in[137]^i_stage_6_comp_in[649];
assign o_stage_6_comp_out[138]=i_stage_6_comp_in[138]^i_stage_6_comp_in[650];
assign o_stage_6_comp_out[139]=i_stage_6_comp_in[139]^i_stage_6_comp_in[651];
assign o_stage_6_comp_out[140]=i_stage_6_comp_in[140]^i_stage_6_comp_in[652];
assign o_stage_6_comp_out[141]=i_stage_6_comp_in[141]^i_stage_6_comp_in[653];
assign o_stage_6_comp_out[142]=i_stage_6_comp_in[142]^i_stage_6_comp_in[654];
assign o_stage_6_comp_out[143]=i_stage_6_comp_in[143]^i_stage_6_comp_in[655];
assign o_stage_6_comp_out[144]=i_stage_6_comp_in[144]^i_stage_6_comp_in[656];
assign o_stage_6_comp_out[145]=i_stage_6_comp_in[145]^i_stage_6_comp_in[657];
assign o_stage_6_comp_out[146]=i_stage_6_comp_in[146]^i_stage_6_comp_in[658];
assign o_stage_6_comp_out[147]=i_stage_6_comp_in[147]^i_stage_6_comp_in[659];
assign o_stage_6_comp_out[148]=i_stage_6_comp_in[148]^i_stage_6_comp_in[660];
assign o_stage_6_comp_out[149]=i_stage_6_comp_in[149]^i_stage_6_comp_in[661];
assign o_stage_6_comp_out[150]=i_stage_6_comp_in[150]^i_stage_6_comp_in[662];
assign o_stage_6_comp_out[151]=i_stage_6_comp_in[151]^i_stage_6_comp_in[663];
assign o_stage_6_comp_out[152]=i_stage_6_comp_in[152]^i_stage_6_comp_in[664];
assign o_stage_6_comp_out[153]=i_stage_6_comp_in[153]^i_stage_6_comp_in[665];
assign o_stage_6_comp_out[154]=i_stage_6_comp_in[154]^i_stage_6_comp_in[666];
assign o_stage_6_comp_out[155]=i_stage_6_comp_in[155]^i_stage_6_comp_in[667];
assign o_stage_6_comp_out[156]=i_stage_6_comp_in[156]^i_stage_6_comp_in[668];
assign o_stage_6_comp_out[157]=i_stage_6_comp_in[157]^i_stage_6_comp_in[669];
assign o_stage_6_comp_out[158]=i_stage_6_comp_in[158]^i_stage_6_comp_in[670];
assign o_stage_6_comp_out[159]=i_stage_6_comp_in[159]^i_stage_6_comp_in[671];
assign o_stage_6_comp_out[160]=i_stage_6_comp_in[160]^i_stage_6_comp_in[672];
assign o_stage_6_comp_out[161]=i_stage_6_comp_in[161]^i_stage_6_comp_in[673];
assign o_stage_6_comp_out[162]=i_stage_6_comp_in[162]^i_stage_6_comp_in[674];
assign o_stage_6_comp_out[163]=i_stage_6_comp_in[163]^i_stage_6_comp_in[675];
assign o_stage_6_comp_out[164]=i_stage_6_comp_in[164]^i_stage_6_comp_in[676];
assign o_stage_6_comp_out[165]=i_stage_6_comp_in[165]^i_stage_6_comp_in[677];
assign o_stage_6_comp_out[166]=i_stage_6_comp_in[166]^i_stage_6_comp_in[678];
assign o_stage_6_comp_out[167]=i_stage_6_comp_in[167]^i_stage_6_comp_in[679];
assign o_stage_6_comp_out[168]=i_stage_6_comp_in[168]^i_stage_6_comp_in[680];
assign o_stage_6_comp_out[169]=i_stage_6_comp_in[169]^i_stage_6_comp_in[681];
assign o_stage_6_comp_out[170]=i_stage_6_comp_in[170]^i_stage_6_comp_in[682];
assign o_stage_6_comp_out[171]=i_stage_6_comp_in[171]^i_stage_6_comp_in[683];
assign o_stage_6_comp_out[172]=i_stage_6_comp_in[172]^i_stage_6_comp_in[684];
assign o_stage_6_comp_out[173]=i_stage_6_comp_in[173]^i_stage_6_comp_in[685];
assign o_stage_6_comp_out[174]=i_stage_6_comp_in[174]^i_stage_6_comp_in[686];
assign o_stage_6_comp_out[175]=i_stage_6_comp_in[175]^i_stage_6_comp_in[687];
assign o_stage_6_comp_out[176]=i_stage_6_comp_in[176]^i_stage_6_comp_in[688];
assign o_stage_6_comp_out[177]=i_stage_6_comp_in[177]^i_stage_6_comp_in[689];
assign o_stage_6_comp_out[178]=i_stage_6_comp_in[178]^i_stage_6_comp_in[690];
assign o_stage_6_comp_out[179]=i_stage_6_comp_in[179]^i_stage_6_comp_in[691];
assign o_stage_6_comp_out[180]=i_stage_6_comp_in[180]^i_stage_6_comp_in[692];
assign o_stage_6_comp_out[181]=i_stage_6_comp_in[181]^i_stage_6_comp_in[693];
assign o_stage_6_comp_out[182]=i_stage_6_comp_in[182]^i_stage_6_comp_in[694];
assign o_stage_6_comp_out[183]=i_stage_6_comp_in[183]^i_stage_6_comp_in[695];
assign o_stage_6_comp_out[184]=i_stage_6_comp_in[184]^i_stage_6_comp_in[696];
assign o_stage_6_comp_out[185]=i_stage_6_comp_in[185]^i_stage_6_comp_in[697];
assign o_stage_6_comp_out[186]=i_stage_6_comp_in[186]^i_stage_6_comp_in[698];
assign o_stage_6_comp_out[187]=i_stage_6_comp_in[187]^i_stage_6_comp_in[699];
assign o_stage_6_comp_out[188]=i_stage_6_comp_in[188]^i_stage_6_comp_in[700];
assign o_stage_6_comp_out[189]=i_stage_6_comp_in[189]^i_stage_6_comp_in[701];
assign o_stage_6_comp_out[190]=i_stage_6_comp_in[190]^i_stage_6_comp_in[702];
assign o_stage_6_comp_out[191]=i_stage_6_comp_in[191]^i_stage_6_comp_in[703];
assign o_stage_6_comp_out[192]=i_stage_6_comp_in[192]^i_stage_6_comp_in[704];
assign o_stage_6_comp_out[193]=i_stage_6_comp_in[193]^i_stage_6_comp_in[705];
assign o_stage_6_comp_out[194]=i_stage_6_comp_in[194]^i_stage_6_comp_in[706];
assign o_stage_6_comp_out[195]=i_stage_6_comp_in[195]^i_stage_6_comp_in[707];
assign o_stage_6_comp_out[196]=i_stage_6_comp_in[196]^i_stage_6_comp_in[708];
assign o_stage_6_comp_out[197]=i_stage_6_comp_in[197]^i_stage_6_comp_in[709];
assign o_stage_6_comp_out[198]=i_stage_6_comp_in[198]^i_stage_6_comp_in[710];
assign o_stage_6_comp_out[199]=i_stage_6_comp_in[199]^i_stage_6_comp_in[711];
assign o_stage_6_comp_out[200]=i_stage_6_comp_in[200]^i_stage_6_comp_in[712];
assign o_stage_6_comp_out[201]=i_stage_6_comp_in[201]^i_stage_6_comp_in[713];
assign o_stage_6_comp_out[202]=i_stage_6_comp_in[202]^i_stage_6_comp_in[714];
assign o_stage_6_comp_out[203]=i_stage_6_comp_in[203]^i_stage_6_comp_in[715];
assign o_stage_6_comp_out[204]=i_stage_6_comp_in[204]^i_stage_6_comp_in[716];
assign o_stage_6_comp_out[205]=i_stage_6_comp_in[205]^i_stage_6_comp_in[717];
assign o_stage_6_comp_out[206]=i_stage_6_comp_in[206]^i_stage_6_comp_in[718];
assign o_stage_6_comp_out[207]=i_stage_6_comp_in[207]^i_stage_6_comp_in[719];
assign o_stage_6_comp_out[208]=i_stage_6_comp_in[208]^i_stage_6_comp_in[720];
assign o_stage_6_comp_out[209]=i_stage_6_comp_in[209]^i_stage_6_comp_in[721];
assign o_stage_6_comp_out[210]=i_stage_6_comp_in[210]^i_stage_6_comp_in[722];
assign o_stage_6_comp_out[211]=i_stage_6_comp_in[211]^i_stage_6_comp_in[723];
assign o_stage_6_comp_out[212]=i_stage_6_comp_in[212]^i_stage_6_comp_in[724];
assign o_stage_6_comp_out[213]=i_stage_6_comp_in[213]^i_stage_6_comp_in[725];
assign o_stage_6_comp_out[214]=i_stage_6_comp_in[214]^i_stage_6_comp_in[726];
assign o_stage_6_comp_out[215]=i_stage_6_comp_in[215]^i_stage_6_comp_in[727];
assign o_stage_6_comp_out[216]=i_stage_6_comp_in[216]^i_stage_6_comp_in[728];
assign o_stage_6_comp_out[217]=i_stage_6_comp_in[217]^i_stage_6_comp_in[729];
assign o_stage_6_comp_out[218]=i_stage_6_comp_in[218]^i_stage_6_comp_in[730];
assign o_stage_6_comp_out[219]=i_stage_6_comp_in[219]^i_stage_6_comp_in[731];
assign o_stage_6_comp_out[220]=i_stage_6_comp_in[220]^i_stage_6_comp_in[732];
assign o_stage_6_comp_out[221]=i_stage_6_comp_in[221]^i_stage_6_comp_in[733];
assign o_stage_6_comp_out[222]=i_stage_6_comp_in[222]^i_stage_6_comp_in[734];
assign o_stage_6_comp_out[223]=i_stage_6_comp_in[223]^i_stage_6_comp_in[735];
assign o_stage_6_comp_out[224]=i_stage_6_comp_in[224]^i_stage_6_comp_in[736];
assign o_stage_6_comp_out[225]=i_stage_6_comp_in[225]^i_stage_6_comp_in[737];
assign o_stage_6_comp_out[226]=i_stage_6_comp_in[226]^i_stage_6_comp_in[738];
assign o_stage_6_comp_out[227]=i_stage_6_comp_in[227]^i_stage_6_comp_in[739];
assign o_stage_6_comp_out[228]=i_stage_6_comp_in[228]^i_stage_6_comp_in[740];
assign o_stage_6_comp_out[229]=i_stage_6_comp_in[229]^i_stage_6_comp_in[741];
assign o_stage_6_comp_out[230]=i_stage_6_comp_in[230]^i_stage_6_comp_in[742];
assign o_stage_6_comp_out[231]=i_stage_6_comp_in[231]^i_stage_6_comp_in[743];
assign o_stage_6_comp_out[232]=i_stage_6_comp_in[232]^i_stage_6_comp_in[744];
assign o_stage_6_comp_out[233]=i_stage_6_comp_in[233]^i_stage_6_comp_in[745];
assign o_stage_6_comp_out[234]=i_stage_6_comp_in[234]^i_stage_6_comp_in[746];
assign o_stage_6_comp_out[235]=i_stage_6_comp_in[235]^i_stage_6_comp_in[747];
assign o_stage_6_comp_out[236]=i_stage_6_comp_in[236]^i_stage_6_comp_in[748];
assign o_stage_6_comp_out[237]=i_stage_6_comp_in[237]^i_stage_6_comp_in[749];
assign o_stage_6_comp_out[238]=i_stage_6_comp_in[238]^i_stage_6_comp_in[750];
assign o_stage_6_comp_out[239]=i_stage_6_comp_in[239]^i_stage_6_comp_in[751];
assign o_stage_6_comp_out[240]=i_stage_6_comp_in[240]^i_stage_6_comp_in[752];
assign o_stage_6_comp_out[241]=i_stage_6_comp_in[241]^i_stage_6_comp_in[753];
assign o_stage_6_comp_out[242]=i_stage_6_comp_in[242]^i_stage_6_comp_in[754];
assign o_stage_6_comp_out[243]=i_stage_6_comp_in[243]^i_stage_6_comp_in[755];
assign o_stage_6_comp_out[244]=i_stage_6_comp_in[244]^i_stage_6_comp_in[756];
assign o_stage_6_comp_out[245]=i_stage_6_comp_in[245]^i_stage_6_comp_in[757];
assign o_stage_6_comp_out[246]=i_stage_6_comp_in[246]^i_stage_6_comp_in[758];
assign o_stage_6_comp_out[247]=i_stage_6_comp_in[247]^i_stage_6_comp_in[759];
assign o_stage_6_comp_out[248]=i_stage_6_comp_in[248]^i_stage_6_comp_in[760];
assign o_stage_6_comp_out[249]=i_stage_6_comp_in[249]^i_stage_6_comp_in[761];
assign o_stage_6_comp_out[250]=i_stage_6_comp_in[250]^i_stage_6_comp_in[762];
assign o_stage_6_comp_out[251]=i_stage_6_comp_in[251]^i_stage_6_comp_in[763];
assign o_stage_6_comp_out[252]=i_stage_6_comp_in[252]^i_stage_6_comp_in[764];
assign o_stage_6_comp_out[253]=i_stage_6_comp_in[253]^i_stage_6_comp_in[765];
assign o_stage_6_comp_out[254]=i_stage_6_comp_in[254]^i_stage_6_comp_in[766];
assign o_stage_6_comp_out[255]=i_stage_6_comp_in[255]^i_stage_6_comp_in[767];
assign o_stage_6_comp_out[256]=i_stage_6_comp_in[256]^i_stage_6_comp_in[768];
assign o_stage_6_comp_out[257]=i_stage_6_comp_in[257]^i_stage_6_comp_in[769];
assign o_stage_6_comp_out[258]=i_stage_6_comp_in[258]^i_stage_6_comp_in[770];
assign o_stage_6_comp_out[259]=i_stage_6_comp_in[259]^i_stage_6_comp_in[771];
assign o_stage_6_comp_out[260]=i_stage_6_comp_in[260]^i_stage_6_comp_in[772];
assign o_stage_6_comp_out[261]=i_stage_6_comp_in[261]^i_stage_6_comp_in[773];
assign o_stage_6_comp_out[262]=i_stage_6_comp_in[262]^i_stage_6_comp_in[774];
assign o_stage_6_comp_out[263]=i_stage_6_comp_in[263]^i_stage_6_comp_in[775];
assign o_stage_6_comp_out[264]=i_stage_6_comp_in[264]^i_stage_6_comp_in[776];
assign o_stage_6_comp_out[265]=i_stage_6_comp_in[265]^i_stage_6_comp_in[777];
assign o_stage_6_comp_out[266]=i_stage_6_comp_in[266]^i_stage_6_comp_in[778];
assign o_stage_6_comp_out[267]=i_stage_6_comp_in[267]^i_stage_6_comp_in[779];
assign o_stage_6_comp_out[268]=i_stage_6_comp_in[268]^i_stage_6_comp_in[780];
assign o_stage_6_comp_out[269]=i_stage_6_comp_in[269]^i_stage_6_comp_in[781];
assign o_stage_6_comp_out[270]=i_stage_6_comp_in[270]^i_stage_6_comp_in[782];
assign o_stage_6_comp_out[271]=i_stage_6_comp_in[271]^i_stage_6_comp_in[783];
assign o_stage_6_comp_out[272]=i_stage_6_comp_in[272]^i_stage_6_comp_in[784];
assign o_stage_6_comp_out[273]=i_stage_6_comp_in[273]^i_stage_6_comp_in[785];
assign o_stage_6_comp_out[274]=i_stage_6_comp_in[274]^i_stage_6_comp_in[786];
assign o_stage_6_comp_out[275]=i_stage_6_comp_in[275]^i_stage_6_comp_in[787];
assign o_stage_6_comp_out[276]=i_stage_6_comp_in[276]^i_stage_6_comp_in[788];
assign o_stage_6_comp_out[277]=i_stage_6_comp_in[277]^i_stage_6_comp_in[789];
assign o_stage_6_comp_out[278]=i_stage_6_comp_in[278]^i_stage_6_comp_in[790];
assign o_stage_6_comp_out[279]=i_stage_6_comp_in[279]^i_stage_6_comp_in[791];
assign o_stage_6_comp_out[280]=i_stage_6_comp_in[280]^i_stage_6_comp_in[792];
assign o_stage_6_comp_out[281]=i_stage_6_comp_in[281]^i_stage_6_comp_in[793];
assign o_stage_6_comp_out[282]=i_stage_6_comp_in[282]^i_stage_6_comp_in[794];
assign o_stage_6_comp_out[283]=i_stage_6_comp_in[283]^i_stage_6_comp_in[795];
assign o_stage_6_comp_out[284]=i_stage_6_comp_in[284]^i_stage_6_comp_in[796];
assign o_stage_6_comp_out[285]=i_stage_6_comp_in[285]^i_stage_6_comp_in[797];
assign o_stage_6_comp_out[286]=i_stage_6_comp_in[286]^i_stage_6_comp_in[798];
assign o_stage_6_comp_out[287]=i_stage_6_comp_in[287]^i_stage_6_comp_in[799];
assign o_stage_6_comp_out[288]=i_stage_6_comp_in[288]^i_stage_6_comp_in[800];
assign o_stage_6_comp_out[289]=i_stage_6_comp_in[289]^i_stage_6_comp_in[801];
assign o_stage_6_comp_out[290]=i_stage_6_comp_in[290]^i_stage_6_comp_in[802];
assign o_stage_6_comp_out[291]=i_stage_6_comp_in[291]^i_stage_6_comp_in[803];
assign o_stage_6_comp_out[292]=i_stage_6_comp_in[292]^i_stage_6_comp_in[804];
assign o_stage_6_comp_out[293]=i_stage_6_comp_in[293]^i_stage_6_comp_in[805];
assign o_stage_6_comp_out[294]=i_stage_6_comp_in[294]^i_stage_6_comp_in[806];
assign o_stage_6_comp_out[295]=i_stage_6_comp_in[295]^i_stage_6_comp_in[807];
assign o_stage_6_comp_out[296]=i_stage_6_comp_in[296]^i_stage_6_comp_in[808];
assign o_stage_6_comp_out[297]=i_stage_6_comp_in[297]^i_stage_6_comp_in[809];
assign o_stage_6_comp_out[298]=i_stage_6_comp_in[298]^i_stage_6_comp_in[810];
assign o_stage_6_comp_out[299]=i_stage_6_comp_in[299]^i_stage_6_comp_in[811];
assign o_stage_6_comp_out[300]=i_stage_6_comp_in[300]^i_stage_6_comp_in[812];
assign o_stage_6_comp_out[301]=i_stage_6_comp_in[301]^i_stage_6_comp_in[813];
assign o_stage_6_comp_out[302]=i_stage_6_comp_in[302]^i_stage_6_comp_in[814];
assign o_stage_6_comp_out[303]=i_stage_6_comp_in[303]^i_stage_6_comp_in[815];
assign o_stage_6_comp_out[304]=i_stage_6_comp_in[304]^i_stage_6_comp_in[816];
assign o_stage_6_comp_out[305]=i_stage_6_comp_in[305]^i_stage_6_comp_in[817];
assign o_stage_6_comp_out[306]=i_stage_6_comp_in[306]^i_stage_6_comp_in[818];
assign o_stage_6_comp_out[307]=i_stage_6_comp_in[307]^i_stage_6_comp_in[819];
assign o_stage_6_comp_out[308]=i_stage_6_comp_in[308]^i_stage_6_comp_in[820];
assign o_stage_6_comp_out[309]=i_stage_6_comp_in[309]^i_stage_6_comp_in[821];
assign o_stage_6_comp_out[310]=i_stage_6_comp_in[310]^i_stage_6_comp_in[822];
assign o_stage_6_comp_out[311]=i_stage_6_comp_in[311]^i_stage_6_comp_in[823];
assign o_stage_6_comp_out[312]=i_stage_6_comp_in[312]^i_stage_6_comp_in[824];
assign o_stage_6_comp_out[313]=i_stage_6_comp_in[313]^i_stage_6_comp_in[825];
assign o_stage_6_comp_out[314]=i_stage_6_comp_in[314]^i_stage_6_comp_in[826];
assign o_stage_6_comp_out[315]=i_stage_6_comp_in[315]^i_stage_6_comp_in[827];
assign o_stage_6_comp_out[316]=i_stage_6_comp_in[316]^i_stage_6_comp_in[828];
assign o_stage_6_comp_out[317]=i_stage_6_comp_in[317]^i_stage_6_comp_in[829];
assign o_stage_6_comp_out[318]=i_stage_6_comp_in[318]^i_stage_6_comp_in[830];
assign o_stage_6_comp_out[319]=i_stage_6_comp_in[319]^i_stage_6_comp_in[831];
assign o_stage_6_comp_out[320]=i_stage_6_comp_in[320]^i_stage_6_comp_in[832];
assign o_stage_6_comp_out[321]=i_stage_6_comp_in[321]^i_stage_6_comp_in[833];
assign o_stage_6_comp_out[322]=i_stage_6_comp_in[322]^i_stage_6_comp_in[834];
assign o_stage_6_comp_out[323]=i_stage_6_comp_in[323]^i_stage_6_comp_in[835];
assign o_stage_6_comp_out[324]=i_stage_6_comp_in[324]^i_stage_6_comp_in[836];
assign o_stage_6_comp_out[325]=i_stage_6_comp_in[325]^i_stage_6_comp_in[837];
assign o_stage_6_comp_out[326]=i_stage_6_comp_in[326]^i_stage_6_comp_in[838];
assign o_stage_6_comp_out[327]=i_stage_6_comp_in[327]^i_stage_6_comp_in[839];
assign o_stage_6_comp_out[328]=i_stage_6_comp_in[328]^i_stage_6_comp_in[840];
assign o_stage_6_comp_out[329]=i_stage_6_comp_in[329]^i_stage_6_comp_in[841];
assign o_stage_6_comp_out[330]=i_stage_6_comp_in[330]^i_stage_6_comp_in[842];
assign o_stage_6_comp_out[331]=i_stage_6_comp_in[331]^i_stage_6_comp_in[843];
assign o_stage_6_comp_out[332]=i_stage_6_comp_in[332]^i_stage_6_comp_in[844];
assign o_stage_6_comp_out[333]=i_stage_6_comp_in[333]^i_stage_6_comp_in[845];
assign o_stage_6_comp_out[334]=i_stage_6_comp_in[334]^i_stage_6_comp_in[846];
assign o_stage_6_comp_out[335]=i_stage_6_comp_in[335]^i_stage_6_comp_in[847];
assign o_stage_6_comp_out[336]=i_stage_6_comp_in[336]^i_stage_6_comp_in[848];
assign o_stage_6_comp_out[337]=i_stage_6_comp_in[337]^i_stage_6_comp_in[849];
assign o_stage_6_comp_out[338]=i_stage_6_comp_in[338]^i_stage_6_comp_in[850];
assign o_stage_6_comp_out[339]=i_stage_6_comp_in[339]^i_stage_6_comp_in[851];
assign o_stage_6_comp_out[340]=i_stage_6_comp_in[340]^i_stage_6_comp_in[852];
assign o_stage_6_comp_out[341]=i_stage_6_comp_in[341]^i_stage_6_comp_in[853];
assign o_stage_6_comp_out[342]=i_stage_6_comp_in[342]^i_stage_6_comp_in[854];
assign o_stage_6_comp_out[343]=i_stage_6_comp_in[343]^i_stage_6_comp_in[855];
assign o_stage_6_comp_out[344]=i_stage_6_comp_in[344]^i_stage_6_comp_in[856];
assign o_stage_6_comp_out[345]=i_stage_6_comp_in[345]^i_stage_6_comp_in[857];
assign o_stage_6_comp_out[346]=i_stage_6_comp_in[346]^i_stage_6_comp_in[858];
assign o_stage_6_comp_out[347]=i_stage_6_comp_in[347]^i_stage_6_comp_in[859];
assign o_stage_6_comp_out[348]=i_stage_6_comp_in[348]^i_stage_6_comp_in[860];
assign o_stage_6_comp_out[349]=i_stage_6_comp_in[349]^i_stage_6_comp_in[861];
assign o_stage_6_comp_out[350]=i_stage_6_comp_in[350]^i_stage_6_comp_in[862];
assign o_stage_6_comp_out[351]=i_stage_6_comp_in[351]^i_stage_6_comp_in[863];
assign o_stage_6_comp_out[352]=i_stage_6_comp_in[352]^i_stage_6_comp_in[864];
assign o_stage_6_comp_out[353]=i_stage_6_comp_in[353]^i_stage_6_comp_in[865];
assign o_stage_6_comp_out[354]=i_stage_6_comp_in[354]^i_stage_6_comp_in[866];
assign o_stage_6_comp_out[355]=i_stage_6_comp_in[355]^i_stage_6_comp_in[867];
assign o_stage_6_comp_out[356]=i_stage_6_comp_in[356]^i_stage_6_comp_in[868];
assign o_stage_6_comp_out[357]=i_stage_6_comp_in[357]^i_stage_6_comp_in[869];
assign o_stage_6_comp_out[358]=i_stage_6_comp_in[358]^i_stage_6_comp_in[870];
assign o_stage_6_comp_out[359]=i_stage_6_comp_in[359]^i_stage_6_comp_in[871];
assign o_stage_6_comp_out[360]=i_stage_6_comp_in[360]^i_stage_6_comp_in[872];
assign o_stage_6_comp_out[361]=i_stage_6_comp_in[361]^i_stage_6_comp_in[873];
assign o_stage_6_comp_out[362]=i_stage_6_comp_in[362]^i_stage_6_comp_in[874];
assign o_stage_6_comp_out[363]=i_stage_6_comp_in[363]^i_stage_6_comp_in[875];
assign o_stage_6_comp_out[364]=i_stage_6_comp_in[364]^i_stage_6_comp_in[876];
assign o_stage_6_comp_out[365]=i_stage_6_comp_in[365]^i_stage_6_comp_in[877];
assign o_stage_6_comp_out[366]=i_stage_6_comp_in[366]^i_stage_6_comp_in[878];
assign o_stage_6_comp_out[367]=i_stage_6_comp_in[367]^i_stage_6_comp_in[879];
assign o_stage_6_comp_out[368]=i_stage_6_comp_in[368]^i_stage_6_comp_in[880];
assign o_stage_6_comp_out[369]=i_stage_6_comp_in[369]^i_stage_6_comp_in[881];
assign o_stage_6_comp_out[370]=i_stage_6_comp_in[370]^i_stage_6_comp_in[882];
assign o_stage_6_comp_out[371]=i_stage_6_comp_in[371]^i_stage_6_comp_in[883];
assign o_stage_6_comp_out[372]=i_stage_6_comp_in[372]^i_stage_6_comp_in[884];
assign o_stage_6_comp_out[373]=i_stage_6_comp_in[373]^i_stage_6_comp_in[885];
assign o_stage_6_comp_out[374]=i_stage_6_comp_in[374]^i_stage_6_comp_in[886];
assign o_stage_6_comp_out[375]=i_stage_6_comp_in[375]^i_stage_6_comp_in[887];
assign o_stage_6_comp_out[376]=i_stage_6_comp_in[376]^i_stage_6_comp_in[888];
assign o_stage_6_comp_out[377]=i_stage_6_comp_in[377]^i_stage_6_comp_in[889];
assign o_stage_6_comp_out[378]=i_stage_6_comp_in[378]^i_stage_6_comp_in[890];
assign o_stage_6_comp_out[379]=i_stage_6_comp_in[379]^i_stage_6_comp_in[891];
assign o_stage_6_comp_out[380]=i_stage_6_comp_in[380]^i_stage_6_comp_in[892];
assign o_stage_6_comp_out[381]=i_stage_6_comp_in[381]^i_stage_6_comp_in[893];
assign o_stage_6_comp_out[382]=i_stage_6_comp_in[382]^i_stage_6_comp_in[894];
assign o_stage_6_comp_out[383]=i_stage_6_comp_in[383]^i_stage_6_comp_in[895];
assign o_stage_6_comp_out[384]=i_stage_6_comp_in[384]^i_stage_6_comp_in[896];
assign o_stage_6_comp_out[385]=i_stage_6_comp_in[385]^i_stage_6_comp_in[897];
assign o_stage_6_comp_out[386]=i_stage_6_comp_in[386]^i_stage_6_comp_in[898];
assign o_stage_6_comp_out[387]=i_stage_6_comp_in[387]^i_stage_6_comp_in[899];
assign o_stage_6_comp_out[388]=i_stage_6_comp_in[388]^i_stage_6_comp_in[900];
assign o_stage_6_comp_out[389]=i_stage_6_comp_in[389]^i_stage_6_comp_in[901];
assign o_stage_6_comp_out[390]=i_stage_6_comp_in[390]^i_stage_6_comp_in[902];
assign o_stage_6_comp_out[391]=i_stage_6_comp_in[391]^i_stage_6_comp_in[903];
assign o_stage_6_comp_out[392]=i_stage_6_comp_in[392]^i_stage_6_comp_in[904];
assign o_stage_6_comp_out[393]=i_stage_6_comp_in[393]^i_stage_6_comp_in[905];
assign o_stage_6_comp_out[394]=i_stage_6_comp_in[394]^i_stage_6_comp_in[906];
assign o_stage_6_comp_out[395]=i_stage_6_comp_in[395]^i_stage_6_comp_in[907];
assign o_stage_6_comp_out[396]=i_stage_6_comp_in[396]^i_stage_6_comp_in[908];
assign o_stage_6_comp_out[397]=i_stage_6_comp_in[397]^i_stage_6_comp_in[909];
assign o_stage_6_comp_out[398]=i_stage_6_comp_in[398]^i_stage_6_comp_in[910];
assign o_stage_6_comp_out[399]=i_stage_6_comp_in[399]^i_stage_6_comp_in[911];
assign o_stage_6_comp_out[400]=i_stage_6_comp_in[400]^i_stage_6_comp_in[912];
assign o_stage_6_comp_out[401]=i_stage_6_comp_in[401]^i_stage_6_comp_in[913];
assign o_stage_6_comp_out[402]=i_stage_6_comp_in[402]^i_stage_6_comp_in[914];
assign o_stage_6_comp_out[403]=i_stage_6_comp_in[403]^i_stage_6_comp_in[915];
assign o_stage_6_comp_out[404]=i_stage_6_comp_in[404]^i_stage_6_comp_in[916];
assign o_stage_6_comp_out[405]=i_stage_6_comp_in[405]^i_stage_6_comp_in[917];
assign o_stage_6_comp_out[406]=i_stage_6_comp_in[406]^i_stage_6_comp_in[918];
assign o_stage_6_comp_out[407]=i_stage_6_comp_in[407]^i_stage_6_comp_in[919];
assign o_stage_6_comp_out[408]=i_stage_6_comp_in[408]^i_stage_6_comp_in[920];
assign o_stage_6_comp_out[409]=i_stage_6_comp_in[409]^i_stage_6_comp_in[921];
assign o_stage_6_comp_out[410]=i_stage_6_comp_in[410]^i_stage_6_comp_in[922];
assign o_stage_6_comp_out[411]=i_stage_6_comp_in[411]^i_stage_6_comp_in[923];
assign o_stage_6_comp_out[412]=i_stage_6_comp_in[412]^i_stage_6_comp_in[924];
assign o_stage_6_comp_out[413]=i_stage_6_comp_in[413]^i_stage_6_comp_in[925];
assign o_stage_6_comp_out[414]=i_stage_6_comp_in[414]^i_stage_6_comp_in[926];
assign o_stage_6_comp_out[415]=i_stage_6_comp_in[415]^i_stage_6_comp_in[927];
assign o_stage_6_comp_out[416]=i_stage_6_comp_in[416]^i_stage_6_comp_in[928];
assign o_stage_6_comp_out[417]=i_stage_6_comp_in[417]^i_stage_6_comp_in[929];
assign o_stage_6_comp_out[418]=i_stage_6_comp_in[418]^i_stage_6_comp_in[930];
assign o_stage_6_comp_out[419]=i_stage_6_comp_in[419]^i_stage_6_comp_in[931];
assign o_stage_6_comp_out[420]=i_stage_6_comp_in[420]^i_stage_6_comp_in[932];
assign o_stage_6_comp_out[421]=i_stage_6_comp_in[421]^i_stage_6_comp_in[933];
assign o_stage_6_comp_out[422]=i_stage_6_comp_in[422]^i_stage_6_comp_in[934];
assign o_stage_6_comp_out[423]=i_stage_6_comp_in[423]^i_stage_6_comp_in[935];
assign o_stage_6_comp_out[424]=i_stage_6_comp_in[424]^i_stage_6_comp_in[936];
assign o_stage_6_comp_out[425]=i_stage_6_comp_in[425]^i_stage_6_comp_in[937];
assign o_stage_6_comp_out[426]=i_stage_6_comp_in[426]^i_stage_6_comp_in[938];
assign o_stage_6_comp_out[427]=i_stage_6_comp_in[427]^i_stage_6_comp_in[939];
assign o_stage_6_comp_out[428]=i_stage_6_comp_in[428]^i_stage_6_comp_in[940];
assign o_stage_6_comp_out[429]=i_stage_6_comp_in[429]^i_stage_6_comp_in[941];
assign o_stage_6_comp_out[430]=i_stage_6_comp_in[430]^i_stage_6_comp_in[942];
assign o_stage_6_comp_out[431]=i_stage_6_comp_in[431]^i_stage_6_comp_in[943];
assign o_stage_6_comp_out[432]=i_stage_6_comp_in[432]^i_stage_6_comp_in[944];
assign o_stage_6_comp_out[433]=i_stage_6_comp_in[433]^i_stage_6_comp_in[945];
assign o_stage_6_comp_out[434]=i_stage_6_comp_in[434]^i_stage_6_comp_in[946];
assign o_stage_6_comp_out[435]=i_stage_6_comp_in[435]^i_stage_6_comp_in[947];
assign o_stage_6_comp_out[436]=i_stage_6_comp_in[436]^i_stage_6_comp_in[948];
assign o_stage_6_comp_out[437]=i_stage_6_comp_in[437]^i_stage_6_comp_in[949];
assign o_stage_6_comp_out[438]=i_stage_6_comp_in[438]^i_stage_6_comp_in[950];
assign o_stage_6_comp_out[439]=i_stage_6_comp_in[439]^i_stage_6_comp_in[951];
assign o_stage_6_comp_out[440]=i_stage_6_comp_in[440]^i_stage_6_comp_in[952];
assign o_stage_6_comp_out[441]=i_stage_6_comp_in[441]^i_stage_6_comp_in[953];
assign o_stage_6_comp_out[442]=i_stage_6_comp_in[442]^i_stage_6_comp_in[954];
assign o_stage_6_comp_out[443]=i_stage_6_comp_in[443]^i_stage_6_comp_in[955];
assign o_stage_6_comp_out[444]=i_stage_6_comp_in[444]^i_stage_6_comp_in[956];
assign o_stage_6_comp_out[445]=i_stage_6_comp_in[445]^i_stage_6_comp_in[957];
assign o_stage_6_comp_out[446]=i_stage_6_comp_in[446]^i_stage_6_comp_in[958];
assign o_stage_6_comp_out[447]=i_stage_6_comp_in[447]^i_stage_6_comp_in[959];
assign o_stage_6_comp_out[448]=i_stage_6_comp_in[448]^i_stage_6_comp_in[960];
assign o_stage_6_comp_out[449]=i_stage_6_comp_in[449]^i_stage_6_comp_in[961];
assign o_stage_6_comp_out[450]=i_stage_6_comp_in[450]^i_stage_6_comp_in[962];
assign o_stage_6_comp_out[451]=i_stage_6_comp_in[451]^i_stage_6_comp_in[963];
assign o_stage_6_comp_out[452]=i_stage_6_comp_in[452]^i_stage_6_comp_in[964];
assign o_stage_6_comp_out[453]=i_stage_6_comp_in[453]^i_stage_6_comp_in[965];
assign o_stage_6_comp_out[454]=i_stage_6_comp_in[454]^i_stage_6_comp_in[966];
assign o_stage_6_comp_out[455]=i_stage_6_comp_in[455]^i_stage_6_comp_in[967];
assign o_stage_6_comp_out[456]=i_stage_6_comp_in[456]^i_stage_6_comp_in[968];
assign o_stage_6_comp_out[457]=i_stage_6_comp_in[457]^i_stage_6_comp_in[969];
assign o_stage_6_comp_out[458]=i_stage_6_comp_in[458]^i_stage_6_comp_in[970];
assign o_stage_6_comp_out[459]=i_stage_6_comp_in[459]^i_stage_6_comp_in[971];
assign o_stage_6_comp_out[460]=i_stage_6_comp_in[460]^i_stage_6_comp_in[972];
assign o_stage_6_comp_out[461]=i_stage_6_comp_in[461]^i_stage_6_comp_in[973];
assign o_stage_6_comp_out[462]=i_stage_6_comp_in[462]^i_stage_6_comp_in[974];
assign o_stage_6_comp_out[463]=i_stage_6_comp_in[463]^i_stage_6_comp_in[975];
assign o_stage_6_comp_out[464]=i_stage_6_comp_in[464]^i_stage_6_comp_in[976];
assign o_stage_6_comp_out[465]=i_stage_6_comp_in[465]^i_stage_6_comp_in[977];
assign o_stage_6_comp_out[466]=i_stage_6_comp_in[466]^i_stage_6_comp_in[978];
assign o_stage_6_comp_out[467]=i_stage_6_comp_in[467]^i_stage_6_comp_in[979];
assign o_stage_6_comp_out[468]=i_stage_6_comp_in[468]^i_stage_6_comp_in[980];
assign o_stage_6_comp_out[469]=i_stage_6_comp_in[469]^i_stage_6_comp_in[981];
assign o_stage_6_comp_out[470]=i_stage_6_comp_in[470]^i_stage_6_comp_in[982];
assign o_stage_6_comp_out[471]=i_stage_6_comp_in[471]^i_stage_6_comp_in[983];
assign o_stage_6_comp_out[472]=i_stage_6_comp_in[472]^i_stage_6_comp_in[984];
assign o_stage_6_comp_out[473]=i_stage_6_comp_in[473]^i_stage_6_comp_in[985];
assign o_stage_6_comp_out[474]=i_stage_6_comp_in[474]^i_stage_6_comp_in[986];
assign o_stage_6_comp_out[475]=i_stage_6_comp_in[475]^i_stage_6_comp_in[987];
assign o_stage_6_comp_out[476]=i_stage_6_comp_in[476]^i_stage_6_comp_in[988];
assign o_stage_6_comp_out[477]=i_stage_6_comp_in[477]^i_stage_6_comp_in[989];
assign o_stage_6_comp_out[478]=i_stage_6_comp_in[478]^i_stage_6_comp_in[990];
assign o_stage_6_comp_out[479]=i_stage_6_comp_in[479]^i_stage_6_comp_in[991];
assign o_stage_6_comp_out[480]=i_stage_6_comp_in[480]^i_stage_6_comp_in[992];
assign o_stage_6_comp_out[481]=i_stage_6_comp_in[481]^i_stage_6_comp_in[993];
assign o_stage_6_comp_out[482]=i_stage_6_comp_in[482]^i_stage_6_comp_in[994];
assign o_stage_6_comp_out[483]=i_stage_6_comp_in[483]^i_stage_6_comp_in[995];
assign o_stage_6_comp_out[484]=i_stage_6_comp_in[484]^i_stage_6_comp_in[996];
assign o_stage_6_comp_out[485]=i_stage_6_comp_in[485]^i_stage_6_comp_in[997];
assign o_stage_6_comp_out[486]=i_stage_6_comp_in[486]^i_stage_6_comp_in[998];
assign o_stage_6_comp_out[487]=i_stage_6_comp_in[487]^i_stage_6_comp_in[999];
assign o_stage_6_comp_out[488]=i_stage_6_comp_in[488]^i_stage_6_comp_in[1000];
assign o_stage_6_comp_out[489]=i_stage_6_comp_in[489]^i_stage_6_comp_in[1001];
assign o_stage_6_comp_out[490]=i_stage_6_comp_in[490]^i_stage_6_comp_in[1002];
assign o_stage_6_comp_out[491]=i_stage_6_comp_in[491]^i_stage_6_comp_in[1003];
assign o_stage_6_comp_out[492]=i_stage_6_comp_in[492]^i_stage_6_comp_in[1004];
assign o_stage_6_comp_out[493]=i_stage_6_comp_in[493]^i_stage_6_comp_in[1005];
assign o_stage_6_comp_out[494]=i_stage_6_comp_in[494]^i_stage_6_comp_in[1006];
assign o_stage_6_comp_out[495]=i_stage_6_comp_in[495]^i_stage_6_comp_in[1007];
assign o_stage_6_comp_out[496]=i_stage_6_comp_in[496]^i_stage_6_comp_in[1008];
assign o_stage_6_comp_out[497]=i_stage_6_comp_in[497]^i_stage_6_comp_in[1009];
assign o_stage_6_comp_out[498]=i_stage_6_comp_in[498]^i_stage_6_comp_in[1010];
assign o_stage_6_comp_out[499]=i_stage_6_comp_in[499]^i_stage_6_comp_in[1011];
assign o_stage_6_comp_out[500]=i_stage_6_comp_in[500]^i_stage_6_comp_in[1012];
assign o_stage_6_comp_out[501]=i_stage_6_comp_in[501]^i_stage_6_comp_in[1013];
assign o_stage_6_comp_out[502]=i_stage_6_comp_in[502]^i_stage_6_comp_in[1014];
assign o_stage_6_comp_out[503]=i_stage_6_comp_in[503]^i_stage_6_comp_in[1015];
assign o_stage_6_comp_out[504]=i_stage_6_comp_in[504]^i_stage_6_comp_in[1016];
assign o_stage_6_comp_out[505]=i_stage_6_comp_in[505]^i_stage_6_comp_in[1017];
assign o_stage_6_comp_out[506]=i_stage_6_comp_in[506]^i_stage_6_comp_in[1018];
assign o_stage_6_comp_out[507]=i_stage_6_comp_in[507]^i_stage_6_comp_in[1019];
assign o_stage_6_comp_out[508]=i_stage_6_comp_in[508]^i_stage_6_comp_in[1020];
assign o_stage_6_comp_out[509]=i_stage_6_comp_in[509]^i_stage_6_comp_in[1021];
assign o_stage_6_comp_out[510]=i_stage_6_comp_in[510]^i_stage_6_comp_in[1022];
assign o_stage_6_comp_out[511]=i_stage_6_comp_in[511]^i_stage_6_comp_in[1023];
assign o_stage_6_comp_out[512]=i_stage_6_comp_in[512];
assign o_stage_6_comp_out[513]=i_stage_6_comp_in[513];
assign o_stage_6_comp_out[514]=i_stage_6_comp_in[514];
assign o_stage_6_comp_out[515]=i_stage_6_comp_in[515];
assign o_stage_6_comp_out[516]=i_stage_6_comp_in[516];
assign o_stage_6_comp_out[517]=i_stage_6_comp_in[517];
assign o_stage_6_comp_out[518]=i_stage_6_comp_in[518];
assign o_stage_6_comp_out[519]=i_stage_6_comp_in[519];
assign o_stage_6_comp_out[520]=i_stage_6_comp_in[520];
assign o_stage_6_comp_out[521]=i_stage_6_comp_in[521];
assign o_stage_6_comp_out[522]=i_stage_6_comp_in[522];
assign o_stage_6_comp_out[523]=i_stage_6_comp_in[523];
assign o_stage_6_comp_out[524]=i_stage_6_comp_in[524];
assign o_stage_6_comp_out[525]=i_stage_6_comp_in[525];
assign o_stage_6_comp_out[526]=i_stage_6_comp_in[526];
assign o_stage_6_comp_out[527]=i_stage_6_comp_in[527];
assign o_stage_6_comp_out[528]=i_stage_6_comp_in[528];
assign o_stage_6_comp_out[529]=i_stage_6_comp_in[529];
assign o_stage_6_comp_out[530]=i_stage_6_comp_in[530];
assign o_stage_6_comp_out[531]=i_stage_6_comp_in[531];
assign o_stage_6_comp_out[532]=i_stage_6_comp_in[532];
assign o_stage_6_comp_out[533]=i_stage_6_comp_in[533];
assign o_stage_6_comp_out[534]=i_stage_6_comp_in[534];
assign o_stage_6_comp_out[535]=i_stage_6_comp_in[535];
assign o_stage_6_comp_out[536]=i_stage_6_comp_in[536];
assign o_stage_6_comp_out[537]=i_stage_6_comp_in[537];
assign o_stage_6_comp_out[538]=i_stage_6_comp_in[538];
assign o_stage_6_comp_out[539]=i_stage_6_comp_in[539];
assign o_stage_6_comp_out[540]=i_stage_6_comp_in[540];
assign o_stage_6_comp_out[541]=i_stage_6_comp_in[541];
assign o_stage_6_comp_out[542]=i_stage_6_comp_in[542];
assign o_stage_6_comp_out[543]=i_stage_6_comp_in[543];
assign o_stage_6_comp_out[544]=i_stage_6_comp_in[544];
assign o_stage_6_comp_out[545]=i_stage_6_comp_in[545];
assign o_stage_6_comp_out[546]=i_stage_6_comp_in[546];
assign o_stage_6_comp_out[547]=i_stage_6_comp_in[547];
assign o_stage_6_comp_out[548]=i_stage_6_comp_in[548];
assign o_stage_6_comp_out[549]=i_stage_6_comp_in[549];
assign o_stage_6_comp_out[550]=i_stage_6_comp_in[550];
assign o_stage_6_comp_out[551]=i_stage_6_comp_in[551];
assign o_stage_6_comp_out[552]=i_stage_6_comp_in[552];
assign o_stage_6_comp_out[553]=i_stage_6_comp_in[553];
assign o_stage_6_comp_out[554]=i_stage_6_comp_in[554];
assign o_stage_6_comp_out[555]=i_stage_6_comp_in[555];
assign o_stage_6_comp_out[556]=i_stage_6_comp_in[556];
assign o_stage_6_comp_out[557]=i_stage_6_comp_in[557];
assign o_stage_6_comp_out[558]=i_stage_6_comp_in[558];
assign o_stage_6_comp_out[559]=i_stage_6_comp_in[559];
assign o_stage_6_comp_out[560]=i_stage_6_comp_in[560];
assign o_stage_6_comp_out[561]=i_stage_6_comp_in[561];
assign o_stage_6_comp_out[562]=i_stage_6_comp_in[562];
assign o_stage_6_comp_out[563]=i_stage_6_comp_in[563];
assign o_stage_6_comp_out[564]=i_stage_6_comp_in[564];
assign o_stage_6_comp_out[565]=i_stage_6_comp_in[565];
assign o_stage_6_comp_out[566]=i_stage_6_comp_in[566];
assign o_stage_6_comp_out[567]=i_stage_6_comp_in[567];
assign o_stage_6_comp_out[568]=i_stage_6_comp_in[568];
assign o_stage_6_comp_out[569]=i_stage_6_comp_in[569];
assign o_stage_6_comp_out[570]=i_stage_6_comp_in[570];
assign o_stage_6_comp_out[571]=i_stage_6_comp_in[571];
assign o_stage_6_comp_out[572]=i_stage_6_comp_in[572];
assign o_stage_6_comp_out[573]=i_stage_6_comp_in[573];
assign o_stage_6_comp_out[574]=i_stage_6_comp_in[574];
assign o_stage_6_comp_out[575]=i_stage_6_comp_in[575];
assign o_stage_6_comp_out[576]=i_stage_6_comp_in[576];
assign o_stage_6_comp_out[577]=i_stage_6_comp_in[577];
assign o_stage_6_comp_out[578]=i_stage_6_comp_in[578];
assign o_stage_6_comp_out[579]=i_stage_6_comp_in[579];
assign o_stage_6_comp_out[580]=i_stage_6_comp_in[580];
assign o_stage_6_comp_out[581]=i_stage_6_comp_in[581];
assign o_stage_6_comp_out[582]=i_stage_6_comp_in[582];
assign o_stage_6_comp_out[583]=i_stage_6_comp_in[583];
assign o_stage_6_comp_out[584]=i_stage_6_comp_in[584];
assign o_stage_6_comp_out[585]=i_stage_6_comp_in[585];
assign o_stage_6_comp_out[586]=i_stage_6_comp_in[586];
assign o_stage_6_comp_out[587]=i_stage_6_comp_in[587];
assign o_stage_6_comp_out[588]=i_stage_6_comp_in[588];
assign o_stage_6_comp_out[589]=i_stage_6_comp_in[589];
assign o_stage_6_comp_out[590]=i_stage_6_comp_in[590];
assign o_stage_6_comp_out[591]=i_stage_6_comp_in[591];
assign o_stage_6_comp_out[592]=i_stage_6_comp_in[592];
assign o_stage_6_comp_out[593]=i_stage_6_comp_in[593];
assign o_stage_6_comp_out[594]=i_stage_6_comp_in[594];
assign o_stage_6_comp_out[595]=i_stage_6_comp_in[595];
assign o_stage_6_comp_out[596]=i_stage_6_comp_in[596];
assign o_stage_6_comp_out[597]=i_stage_6_comp_in[597];
assign o_stage_6_comp_out[598]=i_stage_6_comp_in[598];
assign o_stage_6_comp_out[599]=i_stage_6_comp_in[599];
assign o_stage_6_comp_out[600]=i_stage_6_comp_in[600];
assign o_stage_6_comp_out[601]=i_stage_6_comp_in[601];
assign o_stage_6_comp_out[602]=i_stage_6_comp_in[602];
assign o_stage_6_comp_out[603]=i_stage_6_comp_in[603];
assign o_stage_6_comp_out[604]=i_stage_6_comp_in[604];
assign o_stage_6_comp_out[605]=i_stage_6_comp_in[605];
assign o_stage_6_comp_out[606]=i_stage_6_comp_in[606];
assign o_stage_6_comp_out[607]=i_stage_6_comp_in[607];
assign o_stage_6_comp_out[608]=i_stage_6_comp_in[608];
assign o_stage_6_comp_out[609]=i_stage_6_comp_in[609];
assign o_stage_6_comp_out[610]=i_stage_6_comp_in[610];
assign o_stage_6_comp_out[611]=i_stage_6_comp_in[611];
assign o_stage_6_comp_out[612]=i_stage_6_comp_in[612];
assign o_stage_6_comp_out[613]=i_stage_6_comp_in[613];
assign o_stage_6_comp_out[614]=i_stage_6_comp_in[614];
assign o_stage_6_comp_out[615]=i_stage_6_comp_in[615];
assign o_stage_6_comp_out[616]=i_stage_6_comp_in[616];
assign o_stage_6_comp_out[617]=i_stage_6_comp_in[617];
assign o_stage_6_comp_out[618]=i_stage_6_comp_in[618];
assign o_stage_6_comp_out[619]=i_stage_6_comp_in[619];
assign o_stage_6_comp_out[620]=i_stage_6_comp_in[620];
assign o_stage_6_comp_out[621]=i_stage_6_comp_in[621];
assign o_stage_6_comp_out[622]=i_stage_6_comp_in[622];
assign o_stage_6_comp_out[623]=i_stage_6_comp_in[623];
assign o_stage_6_comp_out[624]=i_stage_6_comp_in[624];
assign o_stage_6_comp_out[625]=i_stage_6_comp_in[625];
assign o_stage_6_comp_out[626]=i_stage_6_comp_in[626];
assign o_stage_6_comp_out[627]=i_stage_6_comp_in[627];
assign o_stage_6_comp_out[628]=i_stage_6_comp_in[628];
assign o_stage_6_comp_out[629]=i_stage_6_comp_in[629];
assign o_stage_6_comp_out[630]=i_stage_6_comp_in[630];
assign o_stage_6_comp_out[631]=i_stage_6_comp_in[631];
assign o_stage_6_comp_out[632]=i_stage_6_comp_in[632];
assign o_stage_6_comp_out[633]=i_stage_6_comp_in[633];
assign o_stage_6_comp_out[634]=i_stage_6_comp_in[634];
assign o_stage_6_comp_out[635]=i_stage_6_comp_in[635];
assign o_stage_6_comp_out[636]=i_stage_6_comp_in[636];
assign o_stage_6_comp_out[637]=i_stage_6_comp_in[637];
assign o_stage_6_comp_out[638]=i_stage_6_comp_in[638];
assign o_stage_6_comp_out[639]=i_stage_6_comp_in[639];
assign o_stage_6_comp_out[640]=i_stage_6_comp_in[640];
assign o_stage_6_comp_out[641]=i_stage_6_comp_in[641];
assign o_stage_6_comp_out[642]=i_stage_6_comp_in[642];
assign o_stage_6_comp_out[643]=i_stage_6_comp_in[643];
assign o_stage_6_comp_out[644]=i_stage_6_comp_in[644];
assign o_stage_6_comp_out[645]=i_stage_6_comp_in[645];
assign o_stage_6_comp_out[646]=i_stage_6_comp_in[646];
assign o_stage_6_comp_out[647]=i_stage_6_comp_in[647];
assign o_stage_6_comp_out[648]=i_stage_6_comp_in[648];
assign o_stage_6_comp_out[649]=i_stage_6_comp_in[649];
assign o_stage_6_comp_out[650]=i_stage_6_comp_in[650];
assign o_stage_6_comp_out[651]=i_stage_6_comp_in[651];
assign o_stage_6_comp_out[652]=i_stage_6_comp_in[652];
assign o_stage_6_comp_out[653]=i_stage_6_comp_in[653];
assign o_stage_6_comp_out[654]=i_stage_6_comp_in[654];
assign o_stage_6_comp_out[655]=i_stage_6_comp_in[655];
assign o_stage_6_comp_out[656]=i_stage_6_comp_in[656];
assign o_stage_6_comp_out[657]=i_stage_6_comp_in[657];
assign o_stage_6_comp_out[658]=i_stage_6_comp_in[658];
assign o_stage_6_comp_out[659]=i_stage_6_comp_in[659];
assign o_stage_6_comp_out[660]=i_stage_6_comp_in[660];
assign o_stage_6_comp_out[661]=i_stage_6_comp_in[661];
assign o_stage_6_comp_out[662]=i_stage_6_comp_in[662];
assign o_stage_6_comp_out[663]=i_stage_6_comp_in[663];
assign o_stage_6_comp_out[664]=i_stage_6_comp_in[664];
assign o_stage_6_comp_out[665]=i_stage_6_comp_in[665];
assign o_stage_6_comp_out[666]=i_stage_6_comp_in[666];
assign o_stage_6_comp_out[667]=i_stage_6_comp_in[667];
assign o_stage_6_comp_out[668]=i_stage_6_comp_in[668];
assign o_stage_6_comp_out[669]=i_stage_6_comp_in[669];
assign o_stage_6_comp_out[670]=i_stage_6_comp_in[670];
assign o_stage_6_comp_out[671]=i_stage_6_comp_in[671];
assign o_stage_6_comp_out[672]=i_stage_6_comp_in[672];
assign o_stage_6_comp_out[673]=i_stage_6_comp_in[673];
assign o_stage_6_comp_out[674]=i_stage_6_comp_in[674];
assign o_stage_6_comp_out[675]=i_stage_6_comp_in[675];
assign o_stage_6_comp_out[676]=i_stage_6_comp_in[676];
assign o_stage_6_comp_out[677]=i_stage_6_comp_in[677];
assign o_stage_6_comp_out[678]=i_stage_6_comp_in[678];
assign o_stage_6_comp_out[679]=i_stage_6_comp_in[679];
assign o_stage_6_comp_out[680]=i_stage_6_comp_in[680];
assign o_stage_6_comp_out[681]=i_stage_6_comp_in[681];
assign o_stage_6_comp_out[682]=i_stage_6_comp_in[682];
assign o_stage_6_comp_out[683]=i_stage_6_comp_in[683];
assign o_stage_6_comp_out[684]=i_stage_6_comp_in[684];
assign o_stage_6_comp_out[685]=i_stage_6_comp_in[685];
assign o_stage_6_comp_out[686]=i_stage_6_comp_in[686];
assign o_stage_6_comp_out[687]=i_stage_6_comp_in[687];
assign o_stage_6_comp_out[688]=i_stage_6_comp_in[688];
assign o_stage_6_comp_out[689]=i_stage_6_comp_in[689];
assign o_stage_6_comp_out[690]=i_stage_6_comp_in[690];
assign o_stage_6_comp_out[691]=i_stage_6_comp_in[691];
assign o_stage_6_comp_out[692]=i_stage_6_comp_in[692];
assign o_stage_6_comp_out[693]=i_stage_6_comp_in[693];
assign o_stage_6_comp_out[694]=i_stage_6_comp_in[694];
assign o_stage_6_comp_out[695]=i_stage_6_comp_in[695];
assign o_stage_6_comp_out[696]=i_stage_6_comp_in[696];
assign o_stage_6_comp_out[697]=i_stage_6_comp_in[697];
assign o_stage_6_comp_out[698]=i_stage_6_comp_in[698];
assign o_stage_6_comp_out[699]=i_stage_6_comp_in[699];
assign o_stage_6_comp_out[700]=i_stage_6_comp_in[700];
assign o_stage_6_comp_out[701]=i_stage_6_comp_in[701];
assign o_stage_6_comp_out[702]=i_stage_6_comp_in[702];
assign o_stage_6_comp_out[703]=i_stage_6_comp_in[703];
assign o_stage_6_comp_out[704]=i_stage_6_comp_in[704];
assign o_stage_6_comp_out[705]=i_stage_6_comp_in[705];
assign o_stage_6_comp_out[706]=i_stage_6_comp_in[706];
assign o_stage_6_comp_out[707]=i_stage_6_comp_in[707];
assign o_stage_6_comp_out[708]=i_stage_6_comp_in[708];
assign o_stage_6_comp_out[709]=i_stage_6_comp_in[709];
assign o_stage_6_comp_out[710]=i_stage_6_comp_in[710];
assign o_stage_6_comp_out[711]=i_stage_6_comp_in[711];
assign o_stage_6_comp_out[712]=i_stage_6_comp_in[712];
assign o_stage_6_comp_out[713]=i_stage_6_comp_in[713];
assign o_stage_6_comp_out[714]=i_stage_6_comp_in[714];
assign o_stage_6_comp_out[715]=i_stage_6_comp_in[715];
assign o_stage_6_comp_out[716]=i_stage_6_comp_in[716];
assign o_stage_6_comp_out[717]=i_stage_6_comp_in[717];
assign o_stage_6_comp_out[718]=i_stage_6_comp_in[718];
assign o_stage_6_comp_out[719]=i_stage_6_comp_in[719];
assign o_stage_6_comp_out[720]=i_stage_6_comp_in[720];
assign o_stage_6_comp_out[721]=i_stage_6_comp_in[721];
assign o_stage_6_comp_out[722]=i_stage_6_comp_in[722];
assign o_stage_6_comp_out[723]=i_stage_6_comp_in[723];
assign o_stage_6_comp_out[724]=i_stage_6_comp_in[724];
assign o_stage_6_comp_out[725]=i_stage_6_comp_in[725];
assign o_stage_6_comp_out[726]=i_stage_6_comp_in[726];
assign o_stage_6_comp_out[727]=i_stage_6_comp_in[727];
assign o_stage_6_comp_out[728]=i_stage_6_comp_in[728];
assign o_stage_6_comp_out[729]=i_stage_6_comp_in[729];
assign o_stage_6_comp_out[730]=i_stage_6_comp_in[730];
assign o_stage_6_comp_out[731]=i_stage_6_comp_in[731];
assign o_stage_6_comp_out[732]=i_stage_6_comp_in[732];
assign o_stage_6_comp_out[733]=i_stage_6_comp_in[733];
assign o_stage_6_comp_out[734]=i_stage_6_comp_in[734];
assign o_stage_6_comp_out[735]=i_stage_6_comp_in[735];
assign o_stage_6_comp_out[736]=i_stage_6_comp_in[736];
assign o_stage_6_comp_out[737]=i_stage_6_comp_in[737];
assign o_stage_6_comp_out[738]=i_stage_6_comp_in[738];
assign o_stage_6_comp_out[739]=i_stage_6_comp_in[739];
assign o_stage_6_comp_out[740]=i_stage_6_comp_in[740];
assign o_stage_6_comp_out[741]=i_stage_6_comp_in[741];
assign o_stage_6_comp_out[742]=i_stage_6_comp_in[742];
assign o_stage_6_comp_out[743]=i_stage_6_comp_in[743];
assign o_stage_6_comp_out[744]=i_stage_6_comp_in[744];
assign o_stage_6_comp_out[745]=i_stage_6_comp_in[745];
assign o_stage_6_comp_out[746]=i_stage_6_comp_in[746];
assign o_stage_6_comp_out[747]=i_stage_6_comp_in[747];
assign o_stage_6_comp_out[748]=i_stage_6_comp_in[748];
assign o_stage_6_comp_out[749]=i_stage_6_comp_in[749];
assign o_stage_6_comp_out[750]=i_stage_6_comp_in[750];
assign o_stage_6_comp_out[751]=i_stage_6_comp_in[751];
assign o_stage_6_comp_out[752]=i_stage_6_comp_in[752];
assign o_stage_6_comp_out[753]=i_stage_6_comp_in[753];
assign o_stage_6_comp_out[754]=i_stage_6_comp_in[754];
assign o_stage_6_comp_out[755]=i_stage_6_comp_in[755];
assign o_stage_6_comp_out[756]=i_stage_6_comp_in[756];
assign o_stage_6_comp_out[757]=i_stage_6_comp_in[757];
assign o_stage_6_comp_out[758]=i_stage_6_comp_in[758];
assign o_stage_6_comp_out[759]=i_stage_6_comp_in[759];
assign o_stage_6_comp_out[760]=i_stage_6_comp_in[760];
assign o_stage_6_comp_out[761]=i_stage_6_comp_in[761];
assign o_stage_6_comp_out[762]=i_stage_6_comp_in[762];
assign o_stage_6_comp_out[763]=i_stage_6_comp_in[763];
assign o_stage_6_comp_out[764]=i_stage_6_comp_in[764];
assign o_stage_6_comp_out[765]=i_stage_6_comp_in[765];
assign o_stage_6_comp_out[766]=i_stage_6_comp_in[766];
assign o_stage_6_comp_out[767]=i_stage_6_comp_in[767];
assign o_stage_6_comp_out[768]=i_stage_6_comp_in[768];
assign o_stage_6_comp_out[769]=i_stage_6_comp_in[769];
assign o_stage_6_comp_out[770]=i_stage_6_comp_in[770];
assign o_stage_6_comp_out[771]=i_stage_6_comp_in[771];
assign o_stage_6_comp_out[772]=i_stage_6_comp_in[772];
assign o_stage_6_comp_out[773]=i_stage_6_comp_in[773];
assign o_stage_6_comp_out[774]=i_stage_6_comp_in[774];
assign o_stage_6_comp_out[775]=i_stage_6_comp_in[775];
assign o_stage_6_comp_out[776]=i_stage_6_comp_in[776];
assign o_stage_6_comp_out[777]=i_stage_6_comp_in[777];
assign o_stage_6_comp_out[778]=i_stage_6_comp_in[778];
assign o_stage_6_comp_out[779]=i_stage_6_comp_in[779];
assign o_stage_6_comp_out[780]=i_stage_6_comp_in[780];
assign o_stage_6_comp_out[781]=i_stage_6_comp_in[781];
assign o_stage_6_comp_out[782]=i_stage_6_comp_in[782];
assign o_stage_6_comp_out[783]=i_stage_6_comp_in[783];
assign o_stage_6_comp_out[784]=i_stage_6_comp_in[784];
assign o_stage_6_comp_out[785]=i_stage_6_comp_in[785];
assign o_stage_6_comp_out[786]=i_stage_6_comp_in[786];
assign o_stage_6_comp_out[787]=i_stage_6_comp_in[787];
assign o_stage_6_comp_out[788]=i_stage_6_comp_in[788];
assign o_stage_6_comp_out[789]=i_stage_6_comp_in[789];
assign o_stage_6_comp_out[790]=i_stage_6_comp_in[790];
assign o_stage_6_comp_out[791]=i_stage_6_comp_in[791];
assign o_stage_6_comp_out[792]=i_stage_6_comp_in[792];
assign o_stage_6_comp_out[793]=i_stage_6_comp_in[793];
assign o_stage_6_comp_out[794]=i_stage_6_comp_in[794];
assign o_stage_6_comp_out[795]=i_stage_6_comp_in[795];
assign o_stage_6_comp_out[796]=i_stage_6_comp_in[796];
assign o_stage_6_comp_out[797]=i_stage_6_comp_in[797];
assign o_stage_6_comp_out[798]=i_stage_6_comp_in[798];
assign o_stage_6_comp_out[799]=i_stage_6_comp_in[799];
assign o_stage_6_comp_out[800]=i_stage_6_comp_in[800];
assign o_stage_6_comp_out[801]=i_stage_6_comp_in[801];
assign o_stage_6_comp_out[802]=i_stage_6_comp_in[802];
assign o_stage_6_comp_out[803]=i_stage_6_comp_in[803];
assign o_stage_6_comp_out[804]=i_stage_6_comp_in[804];
assign o_stage_6_comp_out[805]=i_stage_6_comp_in[805];
assign o_stage_6_comp_out[806]=i_stage_6_comp_in[806];
assign o_stage_6_comp_out[807]=i_stage_6_comp_in[807];
assign o_stage_6_comp_out[808]=i_stage_6_comp_in[808];
assign o_stage_6_comp_out[809]=i_stage_6_comp_in[809];
assign o_stage_6_comp_out[810]=i_stage_6_comp_in[810];
assign o_stage_6_comp_out[811]=i_stage_6_comp_in[811];
assign o_stage_6_comp_out[812]=i_stage_6_comp_in[812];
assign o_stage_6_comp_out[813]=i_stage_6_comp_in[813];
assign o_stage_6_comp_out[814]=i_stage_6_comp_in[814];
assign o_stage_6_comp_out[815]=i_stage_6_comp_in[815];
assign o_stage_6_comp_out[816]=i_stage_6_comp_in[816];
assign o_stage_6_comp_out[817]=i_stage_6_comp_in[817];
assign o_stage_6_comp_out[818]=i_stage_6_comp_in[818];
assign o_stage_6_comp_out[819]=i_stage_6_comp_in[819];
assign o_stage_6_comp_out[820]=i_stage_6_comp_in[820];
assign o_stage_6_comp_out[821]=i_stage_6_comp_in[821];
assign o_stage_6_comp_out[822]=i_stage_6_comp_in[822];
assign o_stage_6_comp_out[823]=i_stage_6_comp_in[823];
assign o_stage_6_comp_out[824]=i_stage_6_comp_in[824];
assign o_stage_6_comp_out[825]=i_stage_6_comp_in[825];
assign o_stage_6_comp_out[826]=i_stage_6_comp_in[826];
assign o_stage_6_comp_out[827]=i_stage_6_comp_in[827];
assign o_stage_6_comp_out[828]=i_stage_6_comp_in[828];
assign o_stage_6_comp_out[829]=i_stage_6_comp_in[829];
assign o_stage_6_comp_out[830]=i_stage_6_comp_in[830];
assign o_stage_6_comp_out[831]=i_stage_6_comp_in[831];
assign o_stage_6_comp_out[832]=i_stage_6_comp_in[832];
assign o_stage_6_comp_out[833]=i_stage_6_comp_in[833];
assign o_stage_6_comp_out[834]=i_stage_6_comp_in[834];
assign o_stage_6_comp_out[835]=i_stage_6_comp_in[835];
assign o_stage_6_comp_out[836]=i_stage_6_comp_in[836];
assign o_stage_6_comp_out[837]=i_stage_6_comp_in[837];
assign o_stage_6_comp_out[838]=i_stage_6_comp_in[838];
assign o_stage_6_comp_out[839]=i_stage_6_comp_in[839];
assign o_stage_6_comp_out[840]=i_stage_6_comp_in[840];
assign o_stage_6_comp_out[841]=i_stage_6_comp_in[841];
assign o_stage_6_comp_out[842]=i_stage_6_comp_in[842];
assign o_stage_6_comp_out[843]=i_stage_6_comp_in[843];
assign o_stage_6_comp_out[844]=i_stage_6_comp_in[844];
assign o_stage_6_comp_out[845]=i_stage_6_comp_in[845];
assign o_stage_6_comp_out[846]=i_stage_6_comp_in[846];
assign o_stage_6_comp_out[847]=i_stage_6_comp_in[847];
assign o_stage_6_comp_out[848]=i_stage_6_comp_in[848];
assign o_stage_6_comp_out[849]=i_stage_6_comp_in[849];
assign o_stage_6_comp_out[850]=i_stage_6_comp_in[850];
assign o_stage_6_comp_out[851]=i_stage_6_comp_in[851];
assign o_stage_6_comp_out[852]=i_stage_6_comp_in[852];
assign o_stage_6_comp_out[853]=i_stage_6_comp_in[853];
assign o_stage_6_comp_out[854]=i_stage_6_comp_in[854];
assign o_stage_6_comp_out[855]=i_stage_6_comp_in[855];
assign o_stage_6_comp_out[856]=i_stage_6_comp_in[856];
assign o_stage_6_comp_out[857]=i_stage_6_comp_in[857];
assign o_stage_6_comp_out[858]=i_stage_6_comp_in[858];
assign o_stage_6_comp_out[859]=i_stage_6_comp_in[859];
assign o_stage_6_comp_out[860]=i_stage_6_comp_in[860];
assign o_stage_6_comp_out[861]=i_stage_6_comp_in[861];
assign o_stage_6_comp_out[862]=i_stage_6_comp_in[862];
assign o_stage_6_comp_out[863]=i_stage_6_comp_in[863];
assign o_stage_6_comp_out[864]=i_stage_6_comp_in[864];
assign o_stage_6_comp_out[865]=i_stage_6_comp_in[865];
assign o_stage_6_comp_out[866]=i_stage_6_comp_in[866];
assign o_stage_6_comp_out[867]=i_stage_6_comp_in[867];
assign o_stage_6_comp_out[868]=i_stage_6_comp_in[868];
assign o_stage_6_comp_out[869]=i_stage_6_comp_in[869];
assign o_stage_6_comp_out[870]=i_stage_6_comp_in[870];
assign o_stage_6_comp_out[871]=i_stage_6_comp_in[871];
assign o_stage_6_comp_out[872]=i_stage_6_comp_in[872];
assign o_stage_6_comp_out[873]=i_stage_6_comp_in[873];
assign o_stage_6_comp_out[874]=i_stage_6_comp_in[874];
assign o_stage_6_comp_out[875]=i_stage_6_comp_in[875];
assign o_stage_6_comp_out[876]=i_stage_6_comp_in[876];
assign o_stage_6_comp_out[877]=i_stage_6_comp_in[877];
assign o_stage_6_comp_out[878]=i_stage_6_comp_in[878];
assign o_stage_6_comp_out[879]=i_stage_6_comp_in[879];
assign o_stage_6_comp_out[880]=i_stage_6_comp_in[880];
assign o_stage_6_comp_out[881]=i_stage_6_comp_in[881];
assign o_stage_6_comp_out[882]=i_stage_6_comp_in[882];
assign o_stage_6_comp_out[883]=i_stage_6_comp_in[883];
assign o_stage_6_comp_out[884]=i_stage_6_comp_in[884];
assign o_stage_6_comp_out[885]=i_stage_6_comp_in[885];
assign o_stage_6_comp_out[886]=i_stage_6_comp_in[886];
assign o_stage_6_comp_out[887]=i_stage_6_comp_in[887];
assign o_stage_6_comp_out[888]=i_stage_6_comp_in[888];
assign o_stage_6_comp_out[889]=i_stage_6_comp_in[889];
assign o_stage_6_comp_out[890]=i_stage_6_comp_in[890];
assign o_stage_6_comp_out[891]=i_stage_6_comp_in[891];
assign o_stage_6_comp_out[892]=i_stage_6_comp_in[892];
assign o_stage_6_comp_out[893]=i_stage_6_comp_in[893];
assign o_stage_6_comp_out[894]=i_stage_6_comp_in[894];
assign o_stage_6_comp_out[895]=i_stage_6_comp_in[895];
assign o_stage_6_comp_out[896]=i_stage_6_comp_in[896];
assign o_stage_6_comp_out[897]=i_stage_6_comp_in[897];
assign o_stage_6_comp_out[898]=i_stage_6_comp_in[898];
assign o_stage_6_comp_out[899]=i_stage_6_comp_in[899];
assign o_stage_6_comp_out[900]=i_stage_6_comp_in[900];
assign o_stage_6_comp_out[901]=i_stage_6_comp_in[901];
assign o_stage_6_comp_out[902]=i_stage_6_comp_in[902];
assign o_stage_6_comp_out[903]=i_stage_6_comp_in[903];
assign o_stage_6_comp_out[904]=i_stage_6_comp_in[904];
assign o_stage_6_comp_out[905]=i_stage_6_comp_in[905];
assign o_stage_6_comp_out[906]=i_stage_6_comp_in[906];
assign o_stage_6_comp_out[907]=i_stage_6_comp_in[907];
assign o_stage_6_comp_out[908]=i_stage_6_comp_in[908];
assign o_stage_6_comp_out[909]=i_stage_6_comp_in[909];
assign o_stage_6_comp_out[910]=i_stage_6_comp_in[910];
assign o_stage_6_comp_out[911]=i_stage_6_comp_in[911];
assign o_stage_6_comp_out[912]=i_stage_6_comp_in[912];
assign o_stage_6_comp_out[913]=i_stage_6_comp_in[913];
assign o_stage_6_comp_out[914]=i_stage_6_comp_in[914];
assign o_stage_6_comp_out[915]=i_stage_6_comp_in[915];
assign o_stage_6_comp_out[916]=i_stage_6_comp_in[916];
assign o_stage_6_comp_out[917]=i_stage_6_comp_in[917];
assign o_stage_6_comp_out[918]=i_stage_6_comp_in[918];
assign o_stage_6_comp_out[919]=i_stage_6_comp_in[919];
assign o_stage_6_comp_out[920]=i_stage_6_comp_in[920];
assign o_stage_6_comp_out[921]=i_stage_6_comp_in[921];
assign o_stage_6_comp_out[922]=i_stage_6_comp_in[922];
assign o_stage_6_comp_out[923]=i_stage_6_comp_in[923];
assign o_stage_6_comp_out[924]=i_stage_6_comp_in[924];
assign o_stage_6_comp_out[925]=i_stage_6_comp_in[925];
assign o_stage_6_comp_out[926]=i_stage_6_comp_in[926];
assign o_stage_6_comp_out[927]=i_stage_6_comp_in[927];
assign o_stage_6_comp_out[928]=i_stage_6_comp_in[928];
assign o_stage_6_comp_out[929]=i_stage_6_comp_in[929];
assign o_stage_6_comp_out[930]=i_stage_6_comp_in[930];
assign o_stage_6_comp_out[931]=i_stage_6_comp_in[931];
assign o_stage_6_comp_out[932]=i_stage_6_comp_in[932];
assign o_stage_6_comp_out[933]=i_stage_6_comp_in[933];
assign o_stage_6_comp_out[934]=i_stage_6_comp_in[934];
assign o_stage_6_comp_out[935]=i_stage_6_comp_in[935];
assign o_stage_6_comp_out[936]=i_stage_6_comp_in[936];
assign o_stage_6_comp_out[937]=i_stage_6_comp_in[937];
assign o_stage_6_comp_out[938]=i_stage_6_comp_in[938];
assign o_stage_6_comp_out[939]=i_stage_6_comp_in[939];
assign o_stage_6_comp_out[940]=i_stage_6_comp_in[940];
assign o_stage_6_comp_out[941]=i_stage_6_comp_in[941];
assign o_stage_6_comp_out[942]=i_stage_6_comp_in[942];
assign o_stage_6_comp_out[943]=i_stage_6_comp_in[943];
assign o_stage_6_comp_out[944]=i_stage_6_comp_in[944];
assign o_stage_6_comp_out[945]=i_stage_6_comp_in[945];
assign o_stage_6_comp_out[946]=i_stage_6_comp_in[946];
assign o_stage_6_comp_out[947]=i_stage_6_comp_in[947];
assign o_stage_6_comp_out[948]=i_stage_6_comp_in[948];
assign o_stage_6_comp_out[949]=i_stage_6_comp_in[949];
assign o_stage_6_comp_out[950]=i_stage_6_comp_in[950];
assign o_stage_6_comp_out[951]=i_stage_6_comp_in[951];
assign o_stage_6_comp_out[952]=i_stage_6_comp_in[952];
assign o_stage_6_comp_out[953]=i_stage_6_comp_in[953];
assign o_stage_6_comp_out[954]=i_stage_6_comp_in[954];
assign o_stage_6_comp_out[955]=i_stage_6_comp_in[955];
assign o_stage_6_comp_out[956]=i_stage_6_comp_in[956];
assign o_stage_6_comp_out[957]=i_stage_6_comp_in[957];
assign o_stage_6_comp_out[958]=i_stage_6_comp_in[958];
assign o_stage_6_comp_out[959]=i_stage_6_comp_in[959];
assign o_stage_6_comp_out[960]=i_stage_6_comp_in[960];
assign o_stage_6_comp_out[961]=i_stage_6_comp_in[961];
assign o_stage_6_comp_out[962]=i_stage_6_comp_in[962];
assign o_stage_6_comp_out[963]=i_stage_6_comp_in[963];
assign o_stage_6_comp_out[964]=i_stage_6_comp_in[964];
assign o_stage_6_comp_out[965]=i_stage_6_comp_in[965];
assign o_stage_6_comp_out[966]=i_stage_6_comp_in[966];
assign o_stage_6_comp_out[967]=i_stage_6_comp_in[967];
assign o_stage_6_comp_out[968]=i_stage_6_comp_in[968];
assign o_stage_6_comp_out[969]=i_stage_6_comp_in[969];
assign o_stage_6_comp_out[970]=i_stage_6_comp_in[970];
assign o_stage_6_comp_out[971]=i_stage_6_comp_in[971];
assign o_stage_6_comp_out[972]=i_stage_6_comp_in[972];
assign o_stage_6_comp_out[973]=i_stage_6_comp_in[973];
assign o_stage_6_comp_out[974]=i_stage_6_comp_in[974];
assign o_stage_6_comp_out[975]=i_stage_6_comp_in[975];
assign o_stage_6_comp_out[976]=i_stage_6_comp_in[976];
assign o_stage_6_comp_out[977]=i_stage_6_comp_in[977];
assign o_stage_6_comp_out[978]=i_stage_6_comp_in[978];
assign o_stage_6_comp_out[979]=i_stage_6_comp_in[979];
assign o_stage_6_comp_out[980]=i_stage_6_comp_in[980];
assign o_stage_6_comp_out[981]=i_stage_6_comp_in[981];
assign o_stage_6_comp_out[982]=i_stage_6_comp_in[982];
assign o_stage_6_comp_out[983]=i_stage_6_comp_in[983];
assign o_stage_6_comp_out[984]=i_stage_6_comp_in[984];
assign o_stage_6_comp_out[985]=i_stage_6_comp_in[985];
assign o_stage_6_comp_out[986]=i_stage_6_comp_in[986];
assign o_stage_6_comp_out[987]=i_stage_6_comp_in[987];
assign o_stage_6_comp_out[988]=i_stage_6_comp_in[988];
assign o_stage_6_comp_out[989]=i_stage_6_comp_in[989];
assign o_stage_6_comp_out[990]=i_stage_6_comp_in[990];
assign o_stage_6_comp_out[991]=i_stage_6_comp_in[991];
assign o_stage_6_comp_out[992]=i_stage_6_comp_in[992];
assign o_stage_6_comp_out[993]=i_stage_6_comp_in[993];
assign o_stage_6_comp_out[994]=i_stage_6_comp_in[994];
assign o_stage_6_comp_out[995]=i_stage_6_comp_in[995];
assign o_stage_6_comp_out[996]=i_stage_6_comp_in[996];
assign o_stage_6_comp_out[997]=i_stage_6_comp_in[997];
assign o_stage_6_comp_out[998]=i_stage_6_comp_in[998];
assign o_stage_6_comp_out[999]=i_stage_6_comp_in[999];
assign o_stage_6_comp_out[1000]=i_stage_6_comp_in[1000];
assign o_stage_6_comp_out[1001]=i_stage_6_comp_in[1001];
assign o_stage_6_comp_out[1002]=i_stage_6_comp_in[1002];
assign o_stage_6_comp_out[1003]=i_stage_6_comp_in[1003];
assign o_stage_6_comp_out[1004]=i_stage_6_comp_in[1004];
assign o_stage_6_comp_out[1005]=i_stage_6_comp_in[1005];
assign o_stage_6_comp_out[1006]=i_stage_6_comp_in[1006];
assign o_stage_6_comp_out[1007]=i_stage_6_comp_in[1007];
assign o_stage_6_comp_out[1008]=i_stage_6_comp_in[1008];
assign o_stage_6_comp_out[1009]=i_stage_6_comp_in[1009];
assign o_stage_6_comp_out[1010]=i_stage_6_comp_in[1010];
assign o_stage_6_comp_out[1011]=i_stage_6_comp_in[1011];
assign o_stage_6_comp_out[1012]=i_stage_6_comp_in[1012];
assign o_stage_6_comp_out[1013]=i_stage_6_comp_in[1013];
assign o_stage_6_comp_out[1014]=i_stage_6_comp_in[1014];
assign o_stage_6_comp_out[1015]=i_stage_6_comp_in[1015];
assign o_stage_6_comp_out[1016]=i_stage_6_comp_in[1016];
assign o_stage_6_comp_out[1017]=i_stage_6_comp_in[1017];
assign o_stage_6_comp_out[1018]=i_stage_6_comp_in[1018];
assign o_stage_6_comp_out[1019]=i_stage_6_comp_in[1019];
assign o_stage_6_comp_out[1020]=i_stage_6_comp_in[1020];
assign o_stage_6_comp_out[1021]=i_stage_6_comp_in[1021];
assign o_stage_6_comp_out[1022]=i_stage_6_comp_in[1022];
assign o_stage_6_comp_out[1023]=i_stage_6_comp_in[1023];


endmodule

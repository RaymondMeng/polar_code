`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Yankai Wang
// 
// Create Date: 2025/05/10 20:02:30
// Design Name: polar_code
// Module Name: Sorter
// Project Name: polar_code
// Target Devices: zcu106
// Tool Versions: 2023.2
// Description: 
//   排序器，输入2L个权重输出筛选后L个最小权重，顺序从小到大
//   排序算法采用简化冒泡排序算法，利用PM特性：
//   PM_{2l} < PM_{2l+1}
//   PM_{2l} < PM_{2l+2}
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//   
//////////////////////////////////////////////////////////////////////////////////
`include "../defines.v"

module Sorter(
    PM_in,
    PM_out
);

/*******************************************************************************/
/*                              Parameter                                      */
/*******************************************************************************/
parameter PM_WIDTH = 8;

`ifdef LIST_SIZE4
    parameter L = 4;
`elsif LIST_SIZE2
    parameter L = 2;
`endif 
/*******************************************************************************/
/*                              IO Direction                                   */
/*******************************************************************************/
input  [PM_WIDTH*2*L-1:0] PM_in;
output [PM_WIDTH*L-1:0]   PM_out;
/*******************************************************************************/
/*                              Signal Declaration                             */
/*******************************************************************************/
/*******************************************************************************/
/*                              Instance                                       */
/*******************************************************************************/
`ifdef LIST_SIZE4
    Sorter4 #(
        .PM_WIDTH(PM_WIDTH)
    ) Sorter4_inst(
        .PM_in(PM_in),
        .PM_out(PM_out)
    );
`elsif LIST_SIZE2
    Sorter2 #(
        .PM_WIDTH(PM_WIDTH)
    ) Sorter2_inst(
        .PM_in(PM_in),
        .PM_out(PM_out)
    );
`endif 
/*******************************************************************************/
/*                              Logic                                          */
/*******************************************************************************/
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Yankai Wang
// 
// Create Date: 2025/05/10 20:02:30
// Design Name: polar_code
// Module Name: PSC
// Project Name: polar_code
// Target Devices: zcu106
// Tool Versions: 2023.2
// Description: 
//   极化码基本单元，x1 = u1 ^ u0, x0 = u0
//   增加使能信号，为1时异或有效，为0时直接输出
//   这里默认索引0为置信度高的比特
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//////////////////////////////////////////////////////////////////////////////////


module PolarBase(
    sel,
    u1,
    u0,
    x1,
    x0
);
/*******************************************************************************/
/*                              Parameter                                      */
/*******************************************************************************/

/*******************************************************************************/
/*                              IO Direction                                   */
/*******************************************************************************/
input  sel;
input  u0, u1;
output x0, x1;
/*******************************************************************************/
/*                              Signal Declaration                             */
/*******************************************************************************/
/*******************************************************************************/
/*                              Instance                                       */
/*******************************************************************************/
/*******************************************************************************/
/*                              Logic                                          */
/*******************************************************************************/
assign x1 = sel ? u0 ^ u1 : u1;
assign x0 = u0; 
endmodule

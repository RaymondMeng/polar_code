`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Yankai Wang
// 
// Create Date: 2025/05/10 20:02:30
// Design Name: polar_code
// Module Name: CAS
// Project Name: polar_code
// Target Devices: zcu106
// Tool Versions: 2023.2
// Description: 
//   Sorter中的比较与交换单元（Compare And Select, CAS）。功能是比较两个输入，将较小的数放在索引低输出
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//   
//////////////////////////////////////////////////////////////////////////////////


module CAS(
    Din0,
    Din1,
    Dout0,
    Dout1
);
/*******************************************************************************/
/*                              Parameter                                      */
/*******************************************************************************/
parameter PM_WIDTH = 8;
/*******************************************************************************/
/*                              IO Direction                                   */
/*******************************************************************************/
input  [PM_WIDTH-1:0] Din0;
input  [PM_WIDTH-1:0] Din1;
output [PM_WIDTH-1:0] Dout0;
output [PM_WIDTH-1:0] Dout1;
/*******************************************************************************/
/*                              Signal Declaration                             */
/*******************************************************************************/
/*******************************************************************************/
/*                              Instance                                       */
/*******************************************************************************/
/*******************************************************************************/
/*                              Logic                                          */
/*******************************************************************************/
assign Dout0 = Din0 < Din1 ? Din0 : Din1;
assign Dout1 = Din0 < Din1 ? Din1 : Din0;
endmodule
